/**
 * This file is part of the Coyote <https://github.com/fpgasystems/Coyote>
 *
 * MIT Licence
 * Copyright (c) 2021-2025, Systems Group, ETH Zurich
 * All rights reserved.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:

 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.

 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
 */

`timescale 1ns / 1ps

import lynxTypes::*;

module logic_reg_array_static #(
    parameter integer       N_STAGES = 2,
    parameter integer       DATA_BITS = AXI_DATA_BITS
) (
	input  logic 			            aclk,
	input  logic 			            aresetn,

    input  logic [DATA_BITS-1:0]        s_data,
    output logic [DATA_BITS-1:0]        m_data
);

logic [N_STAGES-1:0][DATA_BITS-1:0] data;
assign data[0] = s_data;
assign m_data = data[N_STAGES-1];

always_ff @(posedge aclk) begin
    if(~aresetn) begin
        for(int i = 1; i < N_STAGES; i++) 
            data[i] <= 0;
    end 
    else begin
        for(int i = 1; i < N_STAGES; i++) 
            data[i] <= data[i-1];
    end
end

endmodule