-------------------------------------------------------------------------------
-- MSB-first 512b CRC24, generator 0x328B63
-- ./crcgen -P "x^21 + x^20 + x^17 + x^15 + x^11 + x^9 + x^8 + x^6 + x^5 + x + 1" -B 24 -b 512 -V -L -n crc_512_24_328b63 -D X -C R -o R_n
--
-- Copyright (c) 2022 ETH Zurich.
-- All rights reserved.
--
-- This file is distributed under the terms in the attached LICENSE file.
-- If you do not find this file, copies can be found by writing to:
-- ETH Zurich D-INFK, Stampfenbachstrasse 114, CH-8092 Zurich. Attn: Systems Group
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity crc_512_24_328b63 is
port (
    R   :  in std_logic_vector(23 downto 0);
    X   :  in std_logic_vector(511 downto 0);
    R_n : out std_logic_vector(23 downto 0)
);
end crc_512_24_328b63;

architecture functional of crc_512_24_328b63 is
begin

R_n(0) <= (R(0) xor R(4) xor R(5) xor R(6) xor R(7) xor R(11) xor R(12) xor R(13) xor R(14) xor R(15) xor R(18) xor R(19) xor R(21) xor R(22) xor R(23) xor X(0) xor X(3) xor X(4) xor X(6) xor X(7) xor X(8) xor X(10) xor X(11) xor X(14) xor X(16) xor X(23) xor X(29) xor X(30) xor X(31) xor X(32) xor X(34) xor X(36) xor X(37) xor X(38) xor X(39) xor X(41) xor X(46) xor X(48) xor X(49) xor X(52) xor X(53) xor X(56) xor X(58) xor X(59) xor X(60) xor X(62) xor X(63) xor X(64) xor X(65) xor X(66) xor X(67) xor X(69) xor X(70) xor X(73) xor X(77) xor X(80) xor X(83) xor X(85) xor X(86) xor X(87) xor X(89) xor X(91) xor X(97) xor X(98) xor X(99) xor X(100) xor X(103) xor X(104) xor X(107) xor X(113) xor X(118) xor X(119) xor X(123) xor X(124) xor X(126) xor X(127) xor X(131) xor X(132) xor X(133) xor X(137) xor X(138) xor X(140) xor X(146) xor X(148) xor X(149) xor X(151) xor X(153) xor X(154) xor X(155) xor X(156) xor X(157) xor X(158) xor X(160) xor X(161) xor X(163) xor X(164) xor X(165) xor X(166) xor X(175) xor X(177) xor X(182) xor X(183) xor X(185) xor X(187) xor X(190) xor X(191) xor X(192) xor X(193) xor X(194) xor X(196) xor X(199) xor X(200) xor X(203) xor X(204) xor X(205) xor X(207) xor X(208) xor X(211) xor X(212) xor X(214) xor X(218) xor X(219) xor X(220) xor X(223) xor X(224) xor X(225) xor X(229) xor X(230) xor X(231) xor X(235) xor X(236) xor X(237) xor X(240) xor X(243) xor X(244) xor X(245) xor X(246) xor X(247) xor X(248) xor X(249) xor X(251) xor X(252) xor X(254) xor X(257) xor X(258) xor X(259) xor X(260) xor X(261) xor X(262) xor X(264) xor X(265) xor X(266) xor X(273) xor X(274) xor X(275) xor X(278) xor X(279) xor X(281) xor X(285) xor X(286) xor X(287) xor X(288) xor X(291) xor X(292) xor X(294) xor X(295) xor X(296) xor X(297) xor X(298) xor X(304) xor X(309) xor X(310) xor X(311) xor X(312) xor X(313) xor X(317) xor X(319) xor X(322) xor X(323) xor X(324) xor X(326) xor X(328) xor X(329) xor X(330) xor X(331) xor X(332) xor X(333) xor X(334) xor X(335) xor X(336) xor X(338) xor X(339) xor X(342) xor X(343) xor X(344) xor X(346) xor X(350) xor X(352) xor X(354) xor X(355) xor X(356) xor X(358) xor X(359) xor X(361) xor X(364) xor X(365) xor X(369) xor X(370) xor X(371) xor X(372) xor X(373) xor X(374) xor X(375) xor X(379) xor X(382) xor X(384) xor X(385) xor X(386) xor X(390) xor X(391) xor X(392) xor X(393) xor X(394) xor X(395) xor X(400) xor X(401) xor X(402) xor X(406) xor X(407) xor X(408) xor X(409) xor X(414) xor X(420) xor X(422) xor X(423) xor X(426) xor X(427) xor X(428) xor X(429) xor X(431) xor X(433) xor X(435) xor X(436) xor X(438) xor X(439) xor X(440) xor X(441) xor X(445) xor X(446) xor X(449) xor X(452) xor X(454) xor X(457) xor X(466) xor X(467) xor X(468) xor X(471) xor X(475) xor X(476) xor X(478) xor X(479) xor X(482) xor X(485) xor X(486) xor X(487) xor X(488) xor X(492) xor X(493) xor X(494) xor X(495) xor X(499) xor X(500) xor X(501) xor X(502) xor X(503) xor X(506) xor X(507) xor X(509) xor X(510) xor X(511));
R_n(1) <= (R(1) xor R(4) xor R(8) xor R(11) xor R(16) xor R(18) xor R(20) xor R(21) xor X(0) xor X(1) xor X(3) xor X(5) xor X(6) xor X(9) xor X(10) xor X(12) xor X(14) xor X(15) xor X(16) xor X(17) xor X(23) xor X(24) xor X(29) xor X(33) xor X(34) xor X(35) xor X(36) xor X(40) xor X(41) xor X(42) xor X(46) xor X(47) xor X(48) xor X(50) xor X(52) xor X(54) xor X(56) xor X(57) xor X(58) xor X(61) xor X(62) xor X(68) xor X(69) xor X(71) xor X(73) xor X(74) xor X(77) xor X(78) xor X(80) xor X(81) xor X(83) xor X(84) xor X(85) xor X(88) xor X(89) xor X(90) xor X(91) xor X(92) xor X(97) xor X(101) xor X(103) xor X(105) xor X(107) xor X(108) xor X(113) xor X(114) xor X(118) xor X(120) xor X(123) xor X(125) xor X(126) xor X(128) xor X(131) xor X(134) xor X(137) xor X(139) xor X(140) xor X(141) xor X(146) xor X(147) xor X(148) xor X(150) xor X(151) xor X(152) xor X(153) xor X(159) xor X(160) xor X(162) xor X(163) xor X(167) xor X(175) xor X(176) xor X(177) xor X(178) xor X(182) xor X(184) xor X(185) xor X(186) xor X(187) xor X(188) xor X(190) xor X(195) xor X(196) xor X(197) xor X(199) xor X(201) xor X(203) xor X(206) xor X(207) xor X(209) xor X(211) xor X(213) xor X(214) xor X(215) xor X(218) xor X(221) xor X(223) xor X(226) xor X(229) xor X(232) xor X(235) xor X(238) xor X(240) xor X(241) xor X(243) xor X(250) xor X(251) xor X(253) xor X(254) xor X(255) xor X(257) xor X(263) xor X(264) xor X(267) xor X(273) xor X(276) xor X(278) xor X(280) xor X(281) xor X(282) xor X(285) xor X(289) xor X(291) xor X(293) xor X(294) xor X(299) xor X(304) xor X(305) xor X(309) xor X(314) xor X(317) xor X(318) xor X(319) xor X(320) xor X(322) xor X(325) xor X(326) xor X(327) xor X(328) xor X(337) xor X(338) xor X(340) xor X(342) xor X(345) xor X(346) xor X(347) xor X(350) xor X(351) xor X(352) xor X(353) xor X(354) xor X(357) xor X(358) xor X(360) xor X(361) xor X(362) xor X(364) xor X(366) xor X(369) xor X(376) xor X(379) xor X(380) xor X(382) xor X(383) xor X(384) xor X(387) xor X(390) xor X(396) xor X(400) xor X(403) xor X(406) xor X(410) xor X(414) xor X(415) xor X(420) xor X(421) xor X(422) xor X(424) xor X(426) xor X(430) xor X(431) xor X(432) xor X(433) xor X(434) xor X(435) xor X(437) xor X(438) xor X(442) xor X(445) xor X(447) xor X(449) xor X(450) xor X(452) xor X(453) xor X(454) xor X(455) xor X(457) xor X(458) xor X(466) xor X(469) xor X(471) xor X(472) xor X(475) xor X(477) xor X(478) xor X(480) xor X(482) xor X(483) xor X(485) xor X(489) xor X(492) xor X(496) xor X(499) xor X(504) xor X(506) xor X(508) xor X(509));
R_n(2) <= (R(2) xor R(5) xor R(9) xor R(12) xor R(17) xor R(19) xor R(21) xor R(22) xor X(1) xor X(2) xor X(4) xor X(6) xor X(7) xor X(10) xor X(11) xor X(13) xor X(15) xor X(16) xor X(17) xor X(18) xor X(24) xor X(25) xor X(30) xor X(34) xor X(35) xor X(36) xor X(37) xor X(41) xor X(42) xor X(43) xor X(47) xor X(48) xor X(49) xor X(51) xor X(53) xor X(55) xor X(57) xor X(58) xor X(59) xor X(62) xor X(63) xor X(69) xor X(70) xor X(72) xor X(74) xor X(75) xor X(78) xor X(79) xor X(81) xor X(82) xor X(84) xor X(85) xor X(86) xor X(89) xor X(90) xor X(91) xor X(92) xor X(93) xor X(98) xor X(102) xor X(104) xor X(106) xor X(108) xor X(109) xor X(114) xor X(115) xor X(119) xor X(121) xor X(124) xor X(126) xor X(127) xor X(129) xor X(132) xor X(135) xor X(138) xor X(140) xor X(141) xor X(142) xor X(147) xor X(148) xor X(149) xor X(151) xor X(152) xor X(153) xor X(154) xor X(160) xor X(161) xor X(163) xor X(164) xor X(168) xor X(176) xor X(177) xor X(178) xor X(179) xor X(183) xor X(185) xor X(186) xor X(187) xor X(188) xor X(189) xor X(191) xor X(196) xor X(197) xor X(198) xor X(200) xor X(202) xor X(204) xor X(207) xor X(208) xor X(210) xor X(212) xor X(214) xor X(215) xor X(216) xor X(219) xor X(222) xor X(224) xor X(227) xor X(230) xor X(233) xor X(236) xor X(239) xor X(241) xor X(242) xor X(244) xor X(251) xor X(252) xor X(254) xor X(255) xor X(256) xor X(258) xor X(264) xor X(265) xor X(268) xor X(274) xor X(277) xor X(279) xor X(281) xor X(282) xor X(283) xor X(286) xor X(290) xor X(292) xor X(294) xor X(295) xor X(300) xor X(305) xor X(306) xor X(310) xor X(315) xor X(318) xor X(319) xor X(320) xor X(321) xor X(323) xor X(326) xor X(327) xor X(328) xor X(329) xor X(338) xor X(339) xor X(341) xor X(343) xor X(346) xor X(347) xor X(348) xor X(351) xor X(352) xor X(353) xor X(354) xor X(355) xor X(358) xor X(359) xor X(361) xor X(362) xor X(363) xor X(365) xor X(367) xor X(370) xor X(377) xor X(380) xor X(381) xor X(383) xor X(384) xor X(385) xor X(388) xor X(391) xor X(397) xor X(401) xor X(404) xor X(407) xor X(411) xor X(415) xor X(416) xor X(421) xor X(422) xor X(423) xor X(425) xor X(427) xor X(431) xor X(432) xor X(433) xor X(434) xor X(435) xor X(436) xor X(438) xor X(439) xor X(443) xor X(446) xor X(448) xor X(450) xor X(451) xor X(453) xor X(454) xor X(455) xor X(456) xor X(458) xor X(459) xor X(467) xor X(470) xor X(472) xor X(473) xor X(476) xor X(478) xor X(479) xor X(481) xor X(483) xor X(484) xor X(486) xor X(490) xor X(493) xor X(497) xor X(500) xor X(505) xor X(507) xor X(509) xor X(510));
R_n(3) <= (R(3) xor R(6) xor R(10) xor R(13) xor R(18) xor R(20) xor R(22) xor R(23) xor X(2) xor X(3) xor X(5) xor X(7) xor X(8) xor X(11) xor X(12) xor X(14) xor X(16) xor X(17) xor X(18) xor X(19) xor X(25) xor X(26) xor X(31) xor X(35) xor X(36) xor X(37) xor X(38) xor X(42) xor X(43) xor X(44) xor X(48) xor X(49) xor X(50) xor X(52) xor X(54) xor X(56) xor X(58) xor X(59) xor X(60) xor X(63) xor X(64) xor X(70) xor X(71) xor X(73) xor X(75) xor X(76) xor X(79) xor X(80) xor X(82) xor X(83) xor X(85) xor X(86) xor X(87) xor X(90) xor X(91) xor X(92) xor X(93) xor X(94) xor X(99) xor X(103) xor X(105) xor X(107) xor X(109) xor X(110) xor X(115) xor X(116) xor X(120) xor X(122) xor X(125) xor X(127) xor X(128) xor X(130) xor X(133) xor X(136) xor X(139) xor X(141) xor X(142) xor X(143) xor X(148) xor X(149) xor X(150) xor X(152) xor X(153) xor X(154) xor X(155) xor X(161) xor X(162) xor X(164) xor X(165) xor X(169) xor X(177) xor X(178) xor X(179) xor X(180) xor X(184) xor X(186) xor X(187) xor X(188) xor X(189) xor X(190) xor X(192) xor X(197) xor X(198) xor X(199) xor X(201) xor X(203) xor X(205) xor X(208) xor X(209) xor X(211) xor X(213) xor X(215) xor X(216) xor X(217) xor X(220) xor X(223) xor X(225) xor X(228) xor X(231) xor X(234) xor X(237) xor X(240) xor X(242) xor X(243) xor X(245) xor X(252) xor X(253) xor X(255) xor X(256) xor X(257) xor X(259) xor X(265) xor X(266) xor X(269) xor X(275) xor X(278) xor X(280) xor X(282) xor X(283) xor X(284) xor X(287) xor X(291) xor X(293) xor X(295) xor X(296) xor X(301) xor X(306) xor X(307) xor X(311) xor X(316) xor X(319) xor X(320) xor X(321) xor X(322) xor X(324) xor X(327) xor X(328) xor X(329) xor X(330) xor X(339) xor X(340) xor X(342) xor X(344) xor X(347) xor X(348) xor X(349) xor X(352) xor X(353) xor X(354) xor X(355) xor X(356) xor X(359) xor X(360) xor X(362) xor X(363) xor X(364) xor X(366) xor X(368) xor X(371) xor X(378) xor X(381) xor X(382) xor X(384) xor X(385) xor X(386) xor X(389) xor X(392) xor X(398) xor X(402) xor X(405) xor X(408) xor X(412) xor X(416) xor X(417) xor X(422) xor X(423) xor X(424) xor X(426) xor X(428) xor X(432) xor X(433) xor X(434) xor X(435) xor X(436) xor X(437) xor X(439) xor X(440) xor X(444) xor X(447) xor X(449) xor X(451) xor X(452) xor X(454) xor X(455) xor X(456) xor X(457) xor X(459) xor X(460) xor X(468) xor X(471) xor X(473) xor X(474) xor X(477) xor X(479) xor X(480) xor X(482) xor X(484) xor X(485) xor X(487) xor X(491) xor X(494) xor X(498) xor X(501) xor X(506) xor X(508) xor X(510) xor X(511));
R_n(4) <= (R(0) xor R(4) xor R(7) xor R(11) xor R(14) xor R(19) xor R(21) xor R(23) xor X(3) xor X(4) xor X(6) xor X(8) xor X(9) xor X(12) xor X(13) xor X(15) xor X(17) xor X(18) xor X(19) xor X(20) xor X(26) xor X(27) xor X(32) xor X(36) xor X(37) xor X(38) xor X(39) xor X(43) xor X(44) xor X(45) xor X(49) xor X(50) xor X(51) xor X(53) xor X(55) xor X(57) xor X(59) xor X(60) xor X(61) xor X(64) xor X(65) xor X(71) xor X(72) xor X(74) xor X(76) xor X(77) xor X(80) xor X(81) xor X(83) xor X(84) xor X(86) xor X(87) xor X(88) xor X(91) xor X(92) xor X(93) xor X(94) xor X(95) xor X(100) xor X(104) xor X(106) xor X(108) xor X(110) xor X(111) xor X(116) xor X(117) xor X(121) xor X(123) xor X(126) xor X(128) xor X(129) xor X(131) xor X(134) xor X(137) xor X(140) xor X(142) xor X(143) xor X(144) xor X(149) xor X(150) xor X(151) xor X(153) xor X(154) xor X(155) xor X(156) xor X(162) xor X(163) xor X(165) xor X(166) xor X(170) xor X(178) xor X(179) xor X(180) xor X(181) xor X(185) xor X(187) xor X(188) xor X(189) xor X(190) xor X(191) xor X(193) xor X(198) xor X(199) xor X(200) xor X(202) xor X(204) xor X(206) xor X(209) xor X(210) xor X(212) xor X(214) xor X(216) xor X(217) xor X(218) xor X(221) xor X(224) xor X(226) xor X(229) xor X(232) xor X(235) xor X(238) xor X(241) xor X(243) xor X(244) xor X(246) xor X(253) xor X(254) xor X(256) xor X(257) xor X(258) xor X(260) xor X(266) xor X(267) xor X(270) xor X(276) xor X(279) xor X(281) xor X(283) xor X(284) xor X(285) xor X(288) xor X(292) xor X(294) xor X(296) xor X(297) xor X(302) xor X(307) xor X(308) xor X(312) xor X(317) xor X(320) xor X(321) xor X(322) xor X(323) xor X(325) xor X(328) xor X(329) xor X(330) xor X(331) xor X(340) xor X(341) xor X(343) xor X(345) xor X(348) xor X(349) xor X(350) xor X(353) xor X(354) xor X(355) xor X(356) xor X(357) xor X(360) xor X(361) xor X(363) xor X(364) xor X(365) xor X(367) xor X(369) xor X(372) xor X(379) xor X(382) xor X(383) xor X(385) xor X(386) xor X(387) xor X(390) xor X(393) xor X(399) xor X(403) xor X(406) xor X(409) xor X(413) xor X(417) xor X(418) xor X(423) xor X(424) xor X(425) xor X(427) xor X(429) xor X(433) xor X(434) xor X(435) xor X(436) xor X(437) xor X(438) xor X(440) xor X(441) xor X(445) xor X(448) xor X(450) xor X(452) xor X(453) xor X(455) xor X(456) xor X(457) xor X(458) xor X(460) xor X(461) xor X(469) xor X(472) xor X(474) xor X(475) xor X(478) xor X(480) xor X(481) xor X(483) xor X(485) xor X(486) xor X(488) xor X(492) xor X(495) xor X(499) xor X(502) xor X(507) xor X(509) xor X(511));
R_n(5) <= (R(0) xor R(1) xor R(4) xor R(6) xor R(7) xor R(8) xor R(11) xor R(13) xor R(14) xor R(18) xor R(19) xor R(20) xor R(21) xor R(23) xor X(0) xor X(3) xor X(5) xor X(6) xor X(8) xor X(9) xor X(11) xor X(13) xor X(18) xor X(19) xor X(20) xor X(21) xor X(23) xor X(27) xor X(28) xor X(29) xor X(30) xor X(31) xor X(32) xor X(33) xor X(34) xor X(36) xor X(40) xor X(41) xor X(44) xor X(45) xor X(48) xor X(49) xor X(50) xor X(51) xor X(53) xor X(54) xor X(59) xor X(61) xor X(63) xor X(64) xor X(67) xor X(69) xor X(70) xor X(72) xor X(75) xor X(78) xor X(80) xor X(81) xor X(82) xor X(83) xor X(84) xor X(86) xor X(88) xor X(91) xor X(92) xor X(93) xor X(94) xor X(95) xor X(96) xor X(97) xor X(98) xor X(99) xor X(100) xor X(101) xor X(103) xor X(104) xor X(105) xor X(109) xor X(111) xor X(112) xor X(113) xor X(117) xor X(119) xor X(122) xor X(123) xor X(126) xor X(129) xor X(130) xor X(131) xor X(133) xor X(135) xor X(137) xor X(140) xor X(141) xor X(143) xor X(144) xor X(145) xor X(146) xor X(148) xor X(149) xor X(150) xor X(152) xor X(153) xor X(158) xor X(160) xor X(161) xor X(165) xor X(167) xor X(171) xor X(175) xor X(177) xor X(179) xor X(180) xor X(181) xor X(183) xor X(185) xor X(186) xor X(187) xor X(188) xor X(189) xor X(193) xor X(196) xor X(201) xor X(204) xor X(208) xor X(210) xor X(212) xor X(213) xor X(214) xor X(215) xor X(217) xor X(220) xor X(222) xor X(223) xor X(224) xor X(227) xor X(229) xor X(231) xor X(233) xor X(235) xor X(237) xor X(239) xor X(240) xor X(242) xor X(243) xor X(246) xor X(248) xor X(249) xor X(251) xor X(252) xor X(255) xor X(260) xor X(262) xor X(264) xor X(265) xor X(266) xor X(267) xor X(268) xor X(271) xor X(273) xor X(274) xor X(275) xor X(277) xor X(278) xor X(279) xor X(280) xor X(281) xor X(282) xor X(284) xor X(287) xor X(288) xor X(289) xor X(291) xor X(292) xor X(293) xor X(294) xor X(296) xor X(303) xor X(304) xor X(308) xor X(310) xor X(311) xor X(312) xor X(317) xor X(318) xor X(319) xor X(321) xor X(328) xor X(333) xor X(334) xor X(335) xor X(336) xor X(338) xor X(339) xor X(341) xor X(343) xor X(349) xor X(351) xor X(352) xor X(357) xor X(359) xor X(362) xor X(366) xor X(368) xor X(369) xor X(371) xor X(372) xor X(374) xor X(375) xor X(379) xor X(380) xor X(382) xor X(383) xor X(385) xor X(387) xor X(388) xor X(390) xor X(392) xor X(393) xor X(395) xor X(401) xor X(402) xor X(404) xor X(406) xor X(408) xor X(409) xor X(410) xor X(418) xor X(419) xor X(420) xor X(422) xor X(423) xor X(424) xor X(425) xor X(427) xor X(429) xor X(430) xor X(431) xor X(433) xor X(434) xor X(437) xor X(440) xor X(442) xor X(445) xor X(451) xor X(452) xor X(453) xor X(456) xor X(458) xor X(459) xor X(461) xor X(462) xor X(466) xor X(467) xor X(468) xor X(470) xor X(471) xor X(473) xor X(478) xor X(481) xor X(484) xor X(485) xor X(488) xor X(489) xor X(492) xor X(494) xor X(495) xor X(496) xor X(499) xor X(501) xor X(502) xor X(506) xor X(507) xor X(508) xor X(509) xor X(511));
R_n(6) <= (R(0) xor R(1) xor R(2) xor R(4) xor R(6) xor R(8) xor R(9) xor R(11) xor R(13) xor R(18) xor R(20) xor R(23) xor X(0) xor X(1) xor X(3) xor X(8) xor X(9) xor X(11) xor X(12) xor X(16) xor X(19) xor X(20) xor X(21) xor X(22) xor X(23) xor X(24) xor X(28) xor X(33) xor X(35) xor X(36) xor X(38) xor X(39) xor X(42) xor X(45) xor X(48) xor X(50) xor X(51) xor X(53) xor X(54) xor X(55) xor X(56) xor X(58) xor X(59) xor X(63) xor X(66) xor X(67) xor X(68) xor X(69) xor X(71) xor X(76) xor X(77) xor X(79) xor X(80) xor X(81) xor X(82) xor X(84) xor X(86) xor X(91) xor X(92) xor X(93) xor X(94) xor X(95) xor X(96) xor X(101) xor X(102) xor X(103) xor X(105) xor X(106) xor X(107) xor X(110) xor X(112) xor X(114) xor X(119) xor X(120) xor X(126) xor X(130) xor X(133) xor X(134) xor X(136) xor X(137) xor X(140) xor X(141) xor X(142) xor X(144) xor X(145) xor X(147) xor X(148) xor X(150) xor X(155) xor X(156) xor X(157) xor X(158) xor X(159) xor X(160) xor X(162) xor X(163) xor X(164) xor X(165) xor X(168) xor X(172) xor X(175) xor X(176) xor X(177) xor X(178) xor X(180) xor X(181) xor X(183) xor X(184) xor X(185) xor X(186) xor X(188) xor X(189) xor X(191) xor X(192) xor X(193) xor X(196) xor X(197) xor X(199) xor X(200) xor X(202) xor X(203) xor X(204) xor X(207) xor X(208) xor X(209) xor X(212) xor X(213) xor X(215) xor X(216) xor X(219) xor X(220) xor X(221) xor X(228) xor X(229) xor X(231) xor X(232) xor X(234) xor X(235) xor X(237) xor X(238) xor X(241) xor X(245) xor X(246) xor X(248) xor X(250) xor X(251) xor X(253) xor X(254) xor X(256) xor X(257) xor X(258) xor X(259) xor X(260) xor X(262) xor X(263) xor X(264) xor X(267) xor X(268) xor X(269) xor X(272) xor X(273) xor X(276) xor X(280) xor X(282) xor X(283) xor X(286) xor X(287) xor X(289) xor X(290) xor X(291) xor X(293) xor X(296) xor X(298) xor X(305) xor X(310) xor X(317) xor X(318) xor X(320) xor X(323) xor X(324) xor X(326) xor X(328) xor X(330) xor X(331) xor X(332) xor X(333) xor X(337) xor X(338) xor X(340) xor X(343) xor X(346) xor X(353) xor X(354) xor X(355) xor X(356) xor X(359) xor X(360) xor X(361) xor X(363) xor X(364) xor X(365) xor X(367) xor X(371) xor X(374) xor X(376) xor X(379) xor X(380) xor X(381) xor X(382) xor X(383) xor X(385) xor X(388) xor X(389) xor X(390) xor X(392) xor X(395) xor X(396) xor X(400) xor X(401) xor X(403) xor X(405) xor X(406) xor X(408) xor X(410) xor X(411) xor X(414) xor X(419) xor X(421) xor X(422) xor X(424) xor X(425) xor X(427) xor X(429) xor X(430) xor X(432) xor X(433) xor X(434) xor X(436) xor X(439) xor X(440) xor X(443) xor X(445) xor X(449) xor X(453) xor X(459) xor X(460) xor X(462) xor X(463) xor X(466) xor X(469) xor X(472) xor X(474) xor X(475) xor X(476) xor X(478) xor X(487) xor X(488) xor X(489) xor X(490) xor X(492) xor X(494) xor X(496) xor X(497) xor X(499) xor X(501) xor X(506) xor X(508) xor X(511));
R_n(7) <= (R(0) xor R(1) xor R(2) xor R(3) xor R(5) xor R(7) xor R(9) xor R(10) xor R(12) xor R(14) xor R(19) xor R(21) xor X(1) xor X(2) xor X(4) xor X(9) xor X(10) xor X(12) xor X(13) xor X(17) xor X(20) xor X(21) xor X(22) xor X(23) xor X(24) xor X(25) xor X(29) xor X(34) xor X(36) xor X(37) xor X(39) xor X(40) xor X(43) xor X(46) xor X(49) xor X(51) xor X(52) xor X(54) xor X(55) xor X(56) xor X(57) xor X(59) xor X(60) xor X(64) xor X(67) xor X(68) xor X(69) xor X(70) xor X(72) xor X(77) xor X(78) xor X(80) xor X(81) xor X(82) xor X(83) xor X(85) xor X(87) xor X(92) xor X(93) xor X(94) xor X(95) xor X(96) xor X(97) xor X(102) xor X(103) xor X(104) xor X(106) xor X(107) xor X(108) xor X(111) xor X(113) xor X(115) xor X(120) xor X(121) xor X(127) xor X(131) xor X(134) xor X(135) xor X(137) xor X(138) xor X(141) xor X(142) xor X(143) xor X(145) xor X(146) xor X(148) xor X(149) xor X(151) xor X(156) xor X(157) xor X(158) xor X(159) xor X(160) xor X(161) xor X(163) xor X(164) xor X(165) xor X(166) xor X(169) xor X(173) xor X(176) xor X(177) xor X(178) xor X(179) xor X(181) xor X(182) xor X(184) xor X(185) xor X(186) xor X(187) xor X(189) xor X(190) xor X(192) xor X(193) xor X(194) xor X(197) xor X(198) xor X(200) xor X(201) xor X(203) xor X(204) xor X(205) xor X(208) xor X(209) xor X(210) xor X(213) xor X(214) xor X(216) xor X(217) xor X(220) xor X(221) xor X(222) xor X(229) xor X(230) xor X(232) xor X(233) xor X(235) xor X(236) xor X(238) xor X(239) xor X(242) xor X(246) xor X(247) xor X(249) xor X(251) xor X(252) xor X(254) xor X(255) xor X(257) xor X(258) xor X(259) xor X(260) xor X(261) xor X(263) xor X(264) xor X(265) xor X(268) xor X(269) xor X(270) xor X(273) xor X(274) xor X(277) xor X(281) xor X(283) xor X(284) xor X(287) xor X(288) xor X(290) xor X(291) xor X(292) xor X(294) xor X(297) xor X(299) xor X(306) xor X(311) xor X(318) xor X(319) xor X(321) xor X(324) xor X(325) xor X(327) xor X(329) xor X(331) xor X(332) xor X(333) xor X(334) xor X(338) xor X(339) xor X(341) xor X(344) xor X(347) xor X(354) xor X(355) xor X(356) xor X(357) xor X(360) xor X(361) xor X(362) xor X(364) xor X(365) xor X(366) xor X(368) xor X(372) xor X(375) xor X(377) xor X(380) xor X(381) xor X(382) xor X(383) xor X(384) xor X(386) xor X(389) xor X(390) xor X(391) xor X(393) xor X(396) xor X(397) xor X(401) xor X(402) xor X(404) xor X(406) xor X(407) xor X(409) xor X(411) xor X(412) xor X(415) xor X(420) xor X(422) xor X(423) xor X(425) xor X(426) xor X(428) xor X(430) xor X(431) xor X(433) xor X(434) xor X(435) xor X(437) xor X(440) xor X(441) xor X(444) xor X(446) xor X(450) xor X(454) xor X(460) xor X(461) xor X(463) xor X(464) xor X(467) xor X(470) xor X(473) xor X(475) xor X(476) xor X(477) xor X(479) xor X(488) xor X(489) xor X(490) xor X(491) xor X(493) xor X(495) xor X(497) xor X(498) xor X(500) xor X(502) xor X(507) xor X(509));
R_n(8) <= (R(0) xor R(1) xor R(2) xor R(3) xor R(5) xor R(7) xor R(8) xor R(10) xor R(12) xor R(14) xor R(18) xor R(19) xor R(20) xor R(21) xor R(23) xor X(0) xor X(2) xor X(4) xor X(5) xor X(6) xor X(7) xor X(8) xor X(13) xor X(16) xor X(18) xor X(21) xor X(22) xor X(24) xor X(25) xor X(26) xor X(29) xor X(31) xor X(32) xor X(34) xor X(35) xor X(36) xor X(39) xor X(40) xor X(44) xor X(46) xor X(47) xor X(48) xor X(49) xor X(50) xor X(55) xor X(57) xor X(59) xor X(61) xor X(62) xor X(63) xor X(64) xor X(66) xor X(67) xor X(68) xor X(71) xor X(77) xor X(78) xor X(79) xor X(80) xor X(81) xor X(82) xor X(84) xor X(85) xor X(87) xor X(88) xor X(89) xor X(91) xor X(93) xor X(94) xor X(95) xor X(96) xor X(99) xor X(100) xor X(105) xor X(108) xor X(109) xor X(112) xor X(113) xor X(114) xor X(116) xor X(118) xor X(119) xor X(121) xor X(122) xor X(123) xor X(124) xor X(126) xor X(127) xor X(128) xor X(131) xor X(133) xor X(135) xor X(136) xor X(137) xor X(139) xor X(140) xor X(142) xor X(143) xor X(144) xor X(147) xor X(148) xor X(150) xor X(151) xor X(152) xor X(153) xor X(154) xor X(155) xor X(156) xor X(159) xor X(162) xor X(163) xor X(167) xor X(170) xor X(174) xor X(175) xor X(178) xor X(179) xor X(180) xor X(186) xor X(188) xor X(192) xor X(195) xor X(196) xor X(198) xor X(200) xor X(201) xor X(202) xor X(203) xor X(206) xor X(207) xor X(208) xor X(209) xor X(210) xor X(212) xor X(215) xor X(217) xor X(219) xor X(220) xor X(221) xor X(222) xor X(224) xor X(225) xor X(229) xor X(233) xor X(234) xor X(235) xor X(239) xor X(244) xor X(245) xor X(246) xor X(249) xor X(250) xor X(251) xor X(253) xor X(254) xor X(255) xor X(256) xor X(257) xor X(269) xor X(270) xor X(271) xor X(273) xor X(279) xor X(281) xor X(282) xor X(284) xor X(286) xor X(287) xor X(289) xor X(293) xor X(294) xor X(296) xor X(297) xor X(300) xor X(304) xor X(307) xor X(309) xor X(310) xor X(311) xor X(313) xor X(317) xor X(320) xor X(323) xor X(324) xor X(325) xor X(329) xor X(331) xor X(336) xor X(338) xor X(340) xor X(343) xor X(344) xor X(345) xor X(346) xor X(348) xor X(350) xor X(352) xor X(354) xor X(357) xor X(359) xor X(362) xor X(363) xor X(364) xor X(366) xor X(367) xor X(370) xor X(371) xor X(372) xor X(374) xor X(375) xor X(376) xor X(378) xor X(379) xor X(381) xor X(383) xor X(386) xor X(387) xor X(393) xor X(395) xor X(397) xor X(398) xor X(400) xor X(401) xor X(403) xor X(405) xor X(406) xor X(409) xor X(410) xor X(412) xor X(413) xor X(414) xor X(416) xor X(420) xor X(421) xor X(422) xor X(424) xor X(428) xor X(432) xor X(433) xor X(434) xor X(439) xor X(440) xor X(442) xor X(446) xor X(447) xor X(449) xor X(451) xor X(452) xor X(454) xor X(455) xor X(457) xor X(461) xor X(462) xor X(464) xor X(465) xor X(466) xor X(467) xor X(474) xor X(475) xor X(477) xor X(479) xor X(480) xor X(482) xor X(485) xor X(486) xor X(487) xor X(488) xor X(489) xor X(490) xor X(491) xor X(493) xor X(495) xor X(496) xor X(498) xor X(500) xor X(502) xor X(506) xor X(507) xor X(508) xor X(509) xor X(511));
R_n(9) <= (R(1) xor R(2) xor R(3) xor R(5) xor R(7) xor R(8) xor R(9) xor R(12) xor R(14) xor R(18) xor R(20) xor R(23) xor X(0) xor X(1) xor X(4) xor X(5) xor X(9) xor X(10) xor X(11) xor X(16) xor X(17) xor X(19) xor X(22) xor X(25) xor X(26) xor X(27) xor X(29) xor X(31) xor X(33) xor X(34) xor X(35) xor X(38) xor X(39) xor X(40) xor X(45) xor X(46) xor X(47) xor X(50) xor X(51) xor X(52) xor X(53) xor X(59) xor X(66) xor X(68) xor X(70) xor X(72) xor X(73) xor X(77) xor X(78) xor X(79) xor X(81) xor X(82) xor X(87) xor X(88) xor X(90) xor X(91) xor X(92) xor X(94) xor X(95) xor X(96) xor X(98) xor X(99) xor X(101) xor X(103) xor X(104) xor X(106) xor X(107) xor X(109) xor X(110) xor X(114) xor X(115) xor X(117) xor X(118) xor X(120) xor X(122) xor X(125) xor X(126) xor X(128) xor X(129) xor X(131) xor X(133) xor X(134) xor X(136) xor X(141) xor X(143) xor X(144) xor X(145) xor X(146) xor X(152) xor X(158) xor X(161) xor X(165) xor X(166) xor X(168) xor X(171) xor X(176) xor X(177) xor X(179) xor X(180) xor X(181) xor X(182) xor X(183) xor X(185) xor X(189) xor X(190) xor X(191) xor X(192) xor X(194) xor X(197) xor X(200) xor X(201) xor X(202) xor X(205) xor X(209) xor X(210) xor X(212) xor X(213) xor X(214) xor X(216) xor X(219) xor X(221) xor X(222) xor X(224) xor X(226) xor X(229) xor X(231) xor X(234) xor X(237) xor X(243) xor X(244) xor X(248) xor X(249) xor X(250) xor X(255) xor X(256) xor X(259) xor X(260) xor X(261) xor X(262) xor X(264) xor X(265) xor X(266) xor X(270) xor X(271) xor X(272) xor X(273) xor X(275) xor X(278) xor X(279) xor X(280) xor X(281) xor X(282) xor X(283) xor X(286) xor X(290) xor X(291) xor X(292) xor X(296) xor X(301) xor X(304) xor X(305) xor X(308) xor X(309) xor X(313) xor X(314) xor X(317) xor X(318) xor X(319) xor X(321) xor X(322) xor X(323) xor X(325) xor X(328) xor X(329) xor X(331) xor X(333) xor X(334) xor X(335) xor X(336) xor X(337) xor X(338) xor X(341) xor X(342) xor X(343) xor X(345) xor X(347) xor X(349) xor X(350) xor X(351) xor X(352) xor X(353) xor X(354) xor X(356) xor X(359) xor X(360) xor X(361) xor X(363) xor X(367) xor X(368) xor X(369) xor X(370) xor X(374) xor X(376) xor X(377) xor X(380) xor X(385) xor X(386) xor X(387) xor X(388) xor X(390) xor X(391) xor X(392) xor X(393) xor X(395) xor X(396) xor X(398) xor X(399) xor X(400) xor X(404) xor X(408) xor X(409) xor X(410) xor X(411) xor X(413) xor X(415) xor X(417) xor X(420) xor X(421) xor X(425) xor X(426) xor X(427) xor X(428) xor X(431) xor X(434) xor X(436) xor X(438) xor X(439) xor X(443) xor X(445) xor X(446) xor X(447) xor X(448) xor X(449) xor X(450) xor X(453) xor X(454) xor X(455) xor X(456) xor X(457) xor X(458) xor X(462) xor X(463) xor X(465) xor X(471) xor X(479) xor X(480) xor X(481) xor X(482) xor X(483) xor X(485) xor X(489) xor X(490) xor X(491) xor X(493) xor X(495) xor X(496) xor X(497) xor X(500) xor X(502) xor X(506) xor X(508) xor X(511));
R_n(10) <= (R(2) xor R(3) xor R(4) xor R(6) xor R(8) xor R(9) xor R(10) xor R(13) xor R(15) xor R(19) xor R(21) xor X(1) xor X(2) xor X(5) xor X(6) xor X(10) xor X(11) xor X(12) xor X(17) xor X(18) xor X(20) xor X(23) xor X(26) xor X(27) xor X(28) xor X(30) xor X(32) xor X(34) xor X(35) xor X(36) xor X(39) xor X(40) xor X(41) xor X(46) xor X(47) xor X(48) xor X(51) xor X(52) xor X(53) xor X(54) xor X(60) xor X(67) xor X(69) xor X(71) xor X(73) xor X(74) xor X(78) xor X(79) xor X(80) xor X(82) xor X(83) xor X(88) xor X(89) xor X(91) xor X(92) xor X(93) xor X(95) xor X(96) xor X(97) xor X(99) xor X(100) xor X(102) xor X(104) xor X(105) xor X(107) xor X(108) xor X(110) xor X(111) xor X(115) xor X(116) xor X(118) xor X(119) xor X(121) xor X(123) xor X(126) xor X(127) xor X(129) xor X(130) xor X(132) xor X(134) xor X(135) xor X(137) xor X(142) xor X(144) xor X(145) xor X(146) xor X(147) xor X(153) xor X(159) xor X(162) xor X(166) xor X(167) xor X(169) xor X(172) xor X(177) xor X(178) xor X(180) xor X(181) xor X(182) xor X(183) xor X(184) xor X(186) xor X(190) xor X(191) xor X(192) xor X(193) xor X(195) xor X(198) xor X(201) xor X(202) xor X(203) xor X(206) xor X(210) xor X(211) xor X(213) xor X(214) xor X(215) xor X(217) xor X(220) xor X(222) xor X(223) xor X(225) xor X(227) xor X(230) xor X(232) xor X(235) xor X(238) xor X(244) xor X(245) xor X(249) xor X(250) xor X(251) xor X(256) xor X(257) xor X(260) xor X(261) xor X(262) xor X(263) xor X(265) xor X(266) xor X(267) xor X(271) xor X(272) xor X(273) xor X(274) xor X(276) xor X(279) xor X(280) xor X(281) xor X(282) xor X(283) xor X(284) xor X(287) xor X(291) xor X(292) xor X(293) xor X(297) xor X(302) xor X(305) xor X(306) xor X(309) xor X(310) xor X(314) xor X(315) xor X(318) xor X(319) xor X(320) xor X(322) xor X(323) xor X(324) xor X(326) xor X(329) xor X(330) xor X(332) xor X(334) xor X(335) xor X(336) xor X(337) xor X(338) xor X(339) xor X(342) xor X(343) xor X(344) xor X(346) xor X(348) xor X(350) xor X(351) xor X(352) xor X(353) xor X(354) xor X(355) xor X(357) xor X(360) xor X(361) xor X(362) xor X(364) xor X(368) xor X(369) xor X(370) xor X(371) xor X(375) xor X(377) xor X(378) xor X(381) xor X(386) xor X(387) xor X(388) xor X(389) xor X(391) xor X(392) xor X(393) xor X(394) xor X(396) xor X(397) xor X(399) xor X(400) xor X(401) xor X(405) xor X(409) xor X(410) xor X(411) xor X(412) xor X(414) xor X(416) xor X(418) xor X(421) xor X(422) xor X(426) xor X(427) xor X(428) xor X(429) xor X(432) xor X(435) xor X(437) xor X(439) xor X(440) xor X(444) xor X(446) xor X(447) xor X(448) xor X(449) xor X(450) xor X(451) xor X(454) xor X(455) xor X(456) xor X(457) xor X(458) xor X(459) xor X(463) xor X(464) xor X(466) xor X(472) xor X(480) xor X(481) xor X(482) xor X(483) xor X(484) xor X(486) xor X(490) xor X(491) xor X(492) xor X(494) xor X(496) xor X(497) xor X(498) xor X(501) xor X(503) xor X(507) xor X(509));
R_n(11) <= (R(0) xor R(3) xor R(6) xor R(9) xor R(10) xor R(12) xor R(13) xor R(15) xor R(16) xor R(18) xor R(19) xor R(20) xor R(21) xor R(23) xor X(0) xor X(2) xor X(4) xor X(8) xor X(10) xor X(12) xor X(13) xor X(14) xor X(16) xor X(18) xor X(19) xor X(21) xor X(23) xor X(24) xor X(27) xor X(28) xor X(30) xor X(32) xor X(33) xor X(34) xor X(35) xor X(38) xor X(39) xor X(40) xor X(42) xor X(46) xor X(47) xor X(54) xor X(55) xor X(56) xor X(58) xor X(59) xor X(60) xor X(61) xor X(62) xor X(63) xor X(64) xor X(65) xor X(66) xor X(67) xor X(68) xor X(69) xor X(72) xor X(73) xor X(74) xor X(75) xor X(77) xor X(79) xor X(81) xor X(84) xor X(85) xor X(86) xor X(87) xor X(90) xor X(91) xor X(92) xor X(93) xor X(94) xor X(96) xor X(99) xor X(101) xor X(104) xor X(105) xor X(106) xor X(107) xor X(108) xor X(109) xor X(111) xor X(112) xor X(113) xor X(116) xor X(117) xor X(118) xor X(120) xor X(122) xor X(123) xor X(126) xor X(128) xor X(130) xor X(132) xor X(135) xor X(136) xor X(137) xor X(140) xor X(143) xor X(145) xor X(147) xor X(149) xor X(151) xor X(153) xor X(155) xor X(156) xor X(157) xor X(158) xor X(161) xor X(164) xor X(165) xor X(166) xor X(167) xor X(168) xor X(170) xor X(173) xor X(175) xor X(177) xor X(178) xor X(179) xor X(181) xor X(184) xor X(190) xor X(200) xor X(202) xor X(205) xor X(208) xor X(215) xor X(216) xor X(219) xor X(220) xor X(221) xor X(225) xor X(226) xor X(228) xor X(229) xor X(230) xor X(233) xor X(235) xor X(237) xor X(239) xor X(240) xor X(243) xor X(244) xor X(247) xor X(248) xor X(249) xor X(250) xor X(254) xor X(259) xor X(260) xor X(263) xor X(265) xor X(267) xor X(268) xor X(272) xor X(277) xor X(278) xor X(279) xor X(280) xor X(282) xor X(283) xor X(284) xor X(286) xor X(287) xor X(291) xor X(293) xor X(295) xor X(296) xor X(297) xor X(303) xor X(304) xor X(306) xor X(307) xor X(309) xor X(312) xor X(313) xor X(315) xor X(316) xor X(317) xor X(320) xor X(321) xor X(322) xor X(325) xor X(326) xor X(327) xor X(328) xor X(329) xor X(332) xor X(334) xor X(337) xor X(340) xor X(342) xor X(345) xor X(346) xor X(347) xor X(349) xor X(350) xor X(351) xor X(353) xor X(359) xor X(362) xor X(363) xor X(364) xor X(373) xor X(374) xor X(375) xor X(376) xor X(378) xor X(384) xor X(385) xor X(386) xor X(387) xor X(388) xor X(389) xor X(391) xor X(397) xor X(398) xor X(407) xor X(408) xor X(409) xor X(410) xor X(411) xor X(412) xor X(413) xor X(414) xor X(415) xor X(417) xor X(419) xor X(420) xor X(426) xor X(430) xor X(431) xor X(435) xor X(439) xor X(446) xor X(447) xor X(448) xor X(450) xor X(451) xor X(454) xor X(455) xor X(456) xor X(458) xor X(459) xor X(460) xor X(464) xor X(465) xor X(466) xor X(468) xor X(471) xor X(473) xor X(475) xor X(476) xor X(478) xor X(479) xor X(481) xor X(483) xor X(484) xor X(486) xor X(488) xor X(491) xor X(494) xor X(497) xor X(498) xor X(500) xor X(501) xor X(503) xor X(504) xor X(506) xor X(507) xor X(508) xor X(509) xor X(511));
R_n(12) <= (R(1) xor R(4) xor R(7) xor R(10) xor R(11) xor R(13) xor R(14) xor R(16) xor R(17) xor R(19) xor R(20) xor R(21) xor R(22) xor X(1) xor X(3) xor X(5) xor X(9) xor X(11) xor X(13) xor X(14) xor X(15) xor X(17) xor X(19) xor X(20) xor X(22) xor X(24) xor X(25) xor X(28) xor X(29) xor X(31) xor X(33) xor X(34) xor X(35) xor X(36) xor X(39) xor X(40) xor X(41) xor X(43) xor X(47) xor X(48) xor X(55) xor X(56) xor X(57) xor X(59) xor X(60) xor X(61) xor X(62) xor X(63) xor X(64) xor X(65) xor X(66) xor X(67) xor X(68) xor X(69) xor X(70) xor X(73) xor X(74) xor X(75) xor X(76) xor X(78) xor X(80) xor X(82) xor X(85) xor X(86) xor X(87) xor X(88) xor X(91) xor X(92) xor X(93) xor X(94) xor X(95) xor X(97) xor X(100) xor X(102) xor X(105) xor X(106) xor X(107) xor X(108) xor X(109) xor X(110) xor X(112) xor X(113) xor X(114) xor X(117) xor X(118) xor X(119) xor X(121) xor X(123) xor X(124) xor X(127) xor X(129) xor X(131) xor X(133) xor X(136) xor X(137) xor X(138) xor X(141) xor X(144) xor X(146) xor X(148) xor X(150) xor X(152) xor X(154) xor X(156) xor X(157) xor X(158) xor X(159) xor X(162) xor X(165) xor X(166) xor X(167) xor X(168) xor X(169) xor X(171) xor X(174) xor X(176) xor X(178) xor X(179) xor X(180) xor X(182) xor X(185) xor X(191) xor X(201) xor X(203) xor X(206) xor X(209) xor X(216) xor X(217) xor X(220) xor X(221) xor X(222) xor X(226) xor X(227) xor X(229) xor X(230) xor X(231) xor X(234) xor X(236) xor X(238) xor X(240) xor X(241) xor X(244) xor X(245) xor X(248) xor X(249) xor X(250) xor X(251) xor X(255) xor X(260) xor X(261) xor X(264) xor X(266) xor X(268) xor X(269) xor X(273) xor X(278) xor X(279) xor X(280) xor X(281) xor X(283) xor X(284) xor X(285) xor X(287) xor X(288) xor X(292) xor X(294) xor X(296) xor X(297) xor X(298) xor X(304) xor X(305) xor X(307) xor X(308) xor X(310) xor X(313) xor X(314) xor X(316) xor X(317) xor X(318) xor X(321) xor X(322) xor X(323) xor X(326) xor X(327) xor X(328) xor X(329) xor X(330) xor X(333) xor X(335) xor X(338) xor X(341) xor X(343) xor X(346) xor X(347) xor X(348) xor X(350) xor X(351) xor X(352) xor X(354) xor X(360) xor X(363) xor X(364) xor X(365) xor X(374) xor X(375) xor X(376) xor X(377) xor X(379) xor X(385) xor X(386) xor X(387) xor X(388) xor X(389) xor X(390) xor X(392) xor X(398) xor X(399) xor X(408) xor X(409) xor X(410) xor X(411) xor X(412) xor X(413) xor X(414) xor X(415) xor X(416) xor X(418) xor X(420) xor X(421) xor X(427) xor X(431) xor X(432) xor X(436) xor X(440) xor X(447) xor X(448) xor X(449) xor X(451) xor X(452) xor X(455) xor X(456) xor X(457) xor X(459) xor X(460) xor X(461) xor X(465) xor X(466) xor X(467) xor X(469) xor X(472) xor X(474) xor X(476) xor X(477) xor X(479) xor X(480) xor X(482) xor X(484) xor X(485) xor X(487) xor X(489) xor X(492) xor X(495) xor X(498) xor X(499) xor X(501) xor X(502) xor X(504) xor X(505) xor X(507) xor X(508) xor X(509) xor X(510));
R_n(13) <= (R(0) xor R(2) xor R(5) xor R(8) xor R(11) xor R(12) xor R(14) xor R(15) xor R(17) xor R(18) xor R(20) xor R(21) xor R(22) xor R(23) xor X(2) xor X(4) xor X(6) xor X(10) xor X(12) xor X(14) xor X(15) xor X(16) xor X(18) xor X(20) xor X(21) xor X(23) xor X(25) xor X(26) xor X(29) xor X(30) xor X(32) xor X(34) xor X(35) xor X(36) xor X(37) xor X(40) xor X(41) xor X(42) xor X(44) xor X(48) xor X(49) xor X(56) xor X(57) xor X(58) xor X(60) xor X(61) xor X(62) xor X(63) xor X(64) xor X(65) xor X(66) xor X(67) xor X(68) xor X(69) xor X(70) xor X(71) xor X(74) xor X(75) xor X(76) xor X(77) xor X(79) xor X(81) xor X(83) xor X(86) xor X(87) xor X(88) xor X(89) xor X(92) xor X(93) xor X(94) xor X(95) xor X(96) xor X(98) xor X(101) xor X(103) xor X(106) xor X(107) xor X(108) xor X(109) xor X(110) xor X(111) xor X(113) xor X(114) xor X(115) xor X(118) xor X(119) xor X(120) xor X(122) xor X(124) xor X(125) xor X(128) xor X(130) xor X(132) xor X(134) xor X(137) xor X(138) xor X(139) xor X(142) xor X(145) xor X(147) xor X(149) xor X(151) xor X(153) xor X(155) xor X(157) xor X(158) xor X(159) xor X(160) xor X(163) xor X(166) xor X(167) xor X(168) xor X(169) xor X(170) xor X(172) xor X(175) xor X(177) xor X(179) xor X(180) xor X(181) xor X(183) xor X(186) xor X(192) xor X(202) xor X(204) xor X(207) xor X(210) xor X(217) xor X(218) xor X(221) xor X(222) xor X(223) xor X(227) xor X(228) xor X(230) xor X(231) xor X(232) xor X(235) xor X(237) xor X(239) xor X(241) xor X(242) xor X(245) xor X(246) xor X(249) xor X(250) xor X(251) xor X(252) xor X(256) xor X(261) xor X(262) xor X(265) xor X(267) xor X(269) xor X(270) xor X(274) xor X(279) xor X(280) xor X(281) xor X(282) xor X(284) xor X(285) xor X(286) xor X(288) xor X(289) xor X(293) xor X(295) xor X(297) xor X(298) xor X(299) xor X(305) xor X(306) xor X(308) xor X(309) xor X(311) xor X(314) xor X(315) xor X(317) xor X(318) xor X(319) xor X(322) xor X(323) xor X(324) xor X(327) xor X(328) xor X(329) xor X(330) xor X(331) xor X(334) xor X(336) xor X(339) xor X(342) xor X(344) xor X(347) xor X(348) xor X(349) xor X(351) xor X(352) xor X(353) xor X(355) xor X(361) xor X(364) xor X(365) xor X(366) xor X(375) xor X(376) xor X(377) xor X(378) xor X(380) xor X(386) xor X(387) xor X(388) xor X(389) xor X(390) xor X(391) xor X(393) xor X(399) xor X(400) xor X(409) xor X(410) xor X(411) xor X(412) xor X(413) xor X(414) xor X(415) xor X(416) xor X(417) xor X(419) xor X(421) xor X(422) xor X(428) xor X(432) xor X(433) xor X(437) xor X(441) xor X(448) xor X(449) xor X(450) xor X(452) xor X(453) xor X(456) xor X(457) xor X(458) xor X(460) xor X(461) xor X(462) xor X(466) xor X(467) xor X(468) xor X(470) xor X(473) xor X(475) xor X(477) xor X(478) xor X(480) xor X(481) xor X(483) xor X(485) xor X(486) xor X(488) xor X(490) xor X(493) xor X(496) xor X(499) xor X(500) xor X(502) xor X(503) xor X(505) xor X(506) xor X(508) xor X(509) xor X(510) xor X(511));
R_n(14) <= (R(1) xor R(3) xor R(6) xor R(9) xor R(12) xor R(13) xor R(15) xor R(16) xor R(18) xor R(19) xor R(21) xor R(22) xor R(23) xor X(3) xor X(5) xor X(7) xor X(11) xor X(13) xor X(15) xor X(16) xor X(17) xor X(19) xor X(21) xor X(22) xor X(24) xor X(26) xor X(27) xor X(30) xor X(31) xor X(33) xor X(35) xor X(36) xor X(37) xor X(38) xor X(41) xor X(42) xor X(43) xor X(45) xor X(49) xor X(50) xor X(57) xor X(58) xor X(59) xor X(61) xor X(62) xor X(63) xor X(64) xor X(65) xor X(66) xor X(67) xor X(68) xor X(69) xor X(70) xor X(71) xor X(72) xor X(75) xor X(76) xor X(77) xor X(78) xor X(80) xor X(82) xor X(84) xor X(87) xor X(88) xor X(89) xor X(90) xor X(93) xor X(94) xor X(95) xor X(96) xor X(97) xor X(99) xor X(102) xor X(104) xor X(107) xor X(108) xor X(109) xor X(110) xor X(111) xor X(112) xor X(114) xor X(115) xor X(116) xor X(119) xor X(120) xor X(121) xor X(123) xor X(125) xor X(126) xor X(129) xor X(131) xor X(133) xor X(135) xor X(138) xor X(139) xor X(140) xor X(143) xor X(146) xor X(148) xor X(150) xor X(152) xor X(154) xor X(156) xor X(158) xor X(159) xor X(160) xor X(161) xor X(164) xor X(167) xor X(168) xor X(169) xor X(170) xor X(171) xor X(173) xor X(176) xor X(178) xor X(180) xor X(181) xor X(182) xor X(184) xor X(187) xor X(193) xor X(203) xor X(205) xor X(208) xor X(211) xor X(218) xor X(219) xor X(222) xor X(223) xor X(224) xor X(228) xor X(229) xor X(231) xor X(232) xor X(233) xor X(236) xor X(238) xor X(240) xor X(242) xor X(243) xor X(246) xor X(247) xor X(250) xor X(251) xor X(252) xor X(253) xor X(257) xor X(262) xor X(263) xor X(266) xor X(268) xor X(270) xor X(271) xor X(275) xor X(280) xor X(281) xor X(282) xor X(283) xor X(285) xor X(286) xor X(287) xor X(289) xor X(290) xor X(294) xor X(296) xor X(298) xor X(299) xor X(300) xor X(306) xor X(307) xor X(309) xor X(310) xor X(312) xor X(315) xor X(316) xor X(318) xor X(319) xor X(320) xor X(323) xor X(324) xor X(325) xor X(328) xor X(329) xor X(330) xor X(331) xor X(332) xor X(335) xor X(337) xor X(340) xor X(343) xor X(345) xor X(348) xor X(349) xor X(350) xor X(352) xor X(353) xor X(354) xor X(356) xor X(362) xor X(365) xor X(366) xor X(367) xor X(376) xor X(377) xor X(378) xor X(379) xor X(381) xor X(387) xor X(388) xor X(389) xor X(390) xor X(391) xor X(392) xor X(394) xor X(400) xor X(401) xor X(410) xor X(411) xor X(412) xor X(413) xor X(414) xor X(415) xor X(416) xor X(417) xor X(418) xor X(420) xor X(422) xor X(423) xor X(429) xor X(433) xor X(434) xor X(438) xor X(442) xor X(449) xor X(450) xor X(451) xor X(453) xor X(454) xor X(457) xor X(458) xor X(459) xor X(461) xor X(462) xor X(463) xor X(467) xor X(468) xor X(469) xor X(471) xor X(474) xor X(476) xor X(478) xor X(479) xor X(481) xor X(482) xor X(484) xor X(486) xor X(487) xor X(489) xor X(491) xor X(494) xor X(497) xor X(500) xor X(501) xor X(503) xor X(504) xor X(506) xor X(507) xor X(509) xor X(510) xor X(511));
R_n(15) <= (R(2) xor R(5) xor R(6) xor R(10) xor R(11) xor R(12) xor R(15) xor R(16) xor R(17) xor R(18) xor R(20) xor R(21) xor X(0) xor X(3) xor X(7) xor X(10) xor X(11) xor X(12) xor X(17) xor X(18) xor X(20) xor X(22) xor X(25) xor X(27) xor X(28) xor X(29) xor X(30) xor X(41) xor X(42) xor X(43) xor X(44) xor X(48) xor X(49) xor X(50) xor X(51) xor X(52) xor X(53) xor X(56) xor X(68) xor X(71) xor X(72) xor X(76) xor X(78) xor X(79) xor X(80) xor X(81) xor X(86) xor X(87) xor X(88) xor X(90) xor X(94) xor X(95) xor X(96) xor X(99) xor X(104) xor X(105) xor X(107) xor X(108) xor X(109) xor X(110) xor X(111) xor X(112) xor X(115) xor X(116) xor X(117) xor X(118) xor X(119) xor X(120) xor X(121) xor X(122) xor X(123) xor X(130) xor X(131) xor X(133) xor X(134) xor X(136) xor X(137) xor X(138) xor X(139) xor X(141) xor X(144) xor X(146) xor X(147) xor X(148) xor X(154) xor X(156) xor X(158) xor X(159) xor X(162) xor X(163) xor X(164) xor X(166) xor X(168) xor X(169) xor X(170) xor X(171) xor X(172) xor X(174) xor X(175) xor X(179) xor X(181) xor X(187) xor X(188) xor X(190) xor X(191) xor X(192) xor X(193) xor X(196) xor X(199) xor X(200) xor X(203) xor X(205) xor X(206) xor X(207) xor X(208) xor X(209) xor X(211) xor X(214) xor X(218) xor X(231) xor X(232) xor X(233) xor X(234) xor X(235) xor X(236) xor X(239) xor X(240) xor X(241) xor X(245) xor X(246) xor X(249) xor X(253) xor X(257) xor X(259) xor X(260) xor X(261) xor X(262) xor X(263) xor X(265) xor X(266) xor X(267) xor X(269) xor X(271) xor X(272) xor X(273) xor X(274) xor X(275) xor X(276) xor X(278) xor X(279) xor X(282) xor X(283) xor X(284) xor X(285) xor X(290) xor X(292) xor X(294) xor X(296) xor X(298) xor X(299) xor X(300) xor X(301) xor X(304) xor X(307) xor X(308) xor X(309) xor X(312) xor X(316) xor X(320) xor X(321) xor X(322) xor X(323) xor X(325) xor X(328) xor X(334) xor X(335) xor X(339) xor X(341) xor X(342) xor X(343) xor X(349) xor X(351) xor X(352) xor X(353) xor X(356) xor X(357) xor X(358) xor X(359) xor X(361) xor X(363) xor X(364) xor X(365) xor X(366) xor X(367) xor X(368) xor X(369) xor X(370) xor X(371) xor X(372) xor X(373) xor X(374) xor X(375) xor X(377) xor X(378) xor X(380) xor X(384) xor X(385) xor X(386) xor X(388) xor X(389) xor X(394) xor X(400) xor X(406) xor X(407) xor X(408) xor X(409) xor X(411) xor X(412) xor X(413) xor X(415) xor X(416) xor X(417) xor X(418) xor X(419) xor X(420) xor X(421) xor X(422) xor X(424) xor X(426) xor X(427) xor X(428) xor X(429) xor X(430) xor X(431) xor X(433) xor X(434) xor X(436) xor X(438) xor X(440) xor X(441) xor X(443) xor X(445) xor X(446) xor X(449) xor X(450) xor X(451) xor X(455) xor X(457) xor X(458) xor X(459) xor X(460) xor X(462) xor X(463) xor X(464) xor X(466) xor X(467) xor X(469) xor X(470) xor X(471) xor X(472) xor X(476) xor X(477) xor X(478) xor X(480) xor X(483) xor X(486) xor X(490) xor X(493) xor X(494) xor X(498) xor X(499) xor X(500) xor X(503) xor X(504) xor X(505) xor X(506) xor X(508) xor X(509));
R_n(16) <= (R(3) xor R(6) xor R(7) xor R(11) xor R(12) xor R(13) xor R(16) xor R(17) xor R(18) xor R(19) xor R(21) xor R(22) xor X(1) xor X(4) xor X(8) xor X(11) xor X(12) xor X(13) xor X(18) xor X(19) xor X(21) xor X(23) xor X(26) xor X(28) xor X(29) xor X(30) xor X(31) xor X(42) xor X(43) xor X(44) xor X(45) xor X(49) xor X(50) xor X(51) xor X(52) xor X(53) xor X(54) xor X(57) xor X(69) xor X(72) xor X(73) xor X(77) xor X(79) xor X(80) xor X(81) xor X(82) xor X(87) xor X(88) xor X(89) xor X(91) xor X(95) xor X(96) xor X(97) xor X(100) xor X(105) xor X(106) xor X(108) xor X(109) xor X(110) xor X(111) xor X(112) xor X(113) xor X(116) xor X(117) xor X(118) xor X(119) xor X(120) xor X(121) xor X(122) xor X(123) xor X(124) xor X(131) xor X(132) xor X(134) xor X(135) xor X(137) xor X(138) xor X(139) xor X(140) xor X(142) xor X(145) xor X(147) xor X(148) xor X(149) xor X(155) xor X(157) xor X(159) xor X(160) xor X(163) xor X(164) xor X(165) xor X(167) xor X(169) xor X(170) xor X(171) xor X(172) xor X(173) xor X(175) xor X(176) xor X(180) xor X(182) xor X(188) xor X(189) xor X(191) xor X(192) xor X(193) xor X(194) xor X(197) xor X(200) xor X(201) xor X(204) xor X(206) xor X(207) xor X(208) xor X(209) xor X(210) xor X(212) xor X(215) xor X(219) xor X(232) xor X(233) xor X(234) xor X(235) xor X(236) xor X(237) xor X(240) xor X(241) xor X(242) xor X(246) xor X(247) xor X(250) xor X(254) xor X(258) xor X(260) xor X(261) xor X(262) xor X(263) xor X(264) xor X(266) xor X(267) xor X(268) xor X(270) xor X(272) xor X(273) xor X(274) xor X(275) xor X(276) xor X(277) xor X(279) xor X(280) xor X(283) xor X(284) xor X(285) xor X(286) xor X(291) xor X(293) xor X(295) xor X(297) xor X(299) xor X(300) xor X(301) xor X(302) xor X(305) xor X(308) xor X(309) xor X(310) xor X(313) xor X(317) xor X(321) xor X(322) xor X(323) xor X(324) xor X(326) xor X(329) xor X(335) xor X(336) xor X(340) xor X(342) xor X(343) xor X(344) xor X(350) xor X(352) xor X(353) xor X(354) xor X(357) xor X(358) xor X(359) xor X(360) xor X(362) xor X(364) xor X(365) xor X(366) xor X(367) xor X(368) xor X(369) xor X(370) xor X(371) xor X(372) xor X(373) xor X(374) xor X(375) xor X(376) xor X(378) xor X(379) xor X(381) xor X(385) xor X(386) xor X(387) xor X(389) xor X(390) xor X(395) xor X(401) xor X(407) xor X(408) xor X(409) xor X(410) xor X(412) xor X(413) xor X(414) xor X(416) xor X(417) xor X(418) xor X(419) xor X(420) xor X(421) xor X(422) xor X(423) xor X(425) xor X(427) xor X(428) xor X(429) xor X(430) xor X(431) xor X(432) xor X(434) xor X(435) xor X(437) xor X(439) xor X(441) xor X(442) xor X(444) xor X(446) xor X(447) xor X(450) xor X(451) xor X(452) xor X(456) xor X(458) xor X(459) xor X(460) xor X(461) xor X(463) xor X(464) xor X(465) xor X(467) xor X(468) xor X(470) xor X(471) xor X(472) xor X(473) xor X(477) xor X(478) xor X(479) xor X(481) xor X(484) xor X(487) xor X(491) xor X(494) xor X(495) xor X(499) xor X(500) xor X(501) xor X(504) xor X(505) xor X(506) xor X(507) xor X(509) xor X(510));
R_n(17) <= (R(5) xor R(6) xor R(8) xor R(11) xor R(15) xor R(17) xor R(20) xor R(21) xor X(0) xor X(2) xor X(3) xor X(4) xor X(5) xor X(6) xor X(7) xor X(8) xor X(9) xor X(10) xor X(11) xor X(12) xor X(13) xor X(16) xor X(19) xor X(20) xor X(22) xor X(23) xor X(24) xor X(27) xor X(34) xor X(36) xor X(37) xor X(38) xor X(39) xor X(41) xor X(43) xor X(44) xor X(45) xor X(48) xor X(49) xor X(50) xor X(51) xor X(54) xor X(55) xor X(56) xor X(59) xor X(60) xor X(62) xor X(63) xor X(64) xor X(65) xor X(66) xor X(67) xor X(69) xor X(74) xor X(77) xor X(78) xor X(81) xor X(82) xor X(85) xor X(86) xor X(87) xor X(88) xor X(90) xor X(91) xor X(92) xor X(96) xor X(99) xor X(100) xor X(101) xor X(103) xor X(104) xor X(106) xor X(109) xor X(110) xor X(111) xor X(112) xor X(114) xor X(117) xor X(120) xor X(121) xor X(122) xor X(125) xor X(126) xor X(127) xor X(131) xor X(135) xor X(136) xor X(137) xor X(139) xor X(141) xor X(143) xor X(150) xor X(151) xor X(153) xor X(154) xor X(155) xor X(157) xor X(163) xor X(168) xor X(170) xor X(171) xor X(172) xor X(173) xor X(174) xor X(175) xor X(176) xor X(181) xor X(182) xor X(185) xor X(187) xor X(189) xor X(191) xor X(195) xor X(196) xor X(198) xor X(199) xor X(200) xor X(201) xor X(202) xor X(203) xor X(204) xor X(209) xor X(210) xor X(212) xor X(213) xor X(214) xor X(216) xor X(218) xor X(219) xor X(223) xor X(224) xor X(225) xor X(229) xor X(230) xor X(231) xor X(233) xor X(234) xor X(238) xor X(240) xor X(241) xor X(242) xor X(244) xor X(245) xor X(246) xor X(249) xor X(252) xor X(254) xor X(255) xor X(257) xor X(258) xor X(260) xor X(263) xor X(266) xor X(267) xor X(268) xor X(269) xor X(271) xor X(276) xor X(277) xor X(279) xor X(280) xor X(284) xor X(288) xor X(291) xor X(295) xor X(297) xor X(300) xor X(301) xor X(302) xor X(303) xor X(304) xor X(306) xor X(312) xor X(313) xor X(314) xor X(317) xor X(318) xor X(319) xor X(325) xor X(326) xor X(327) xor X(328) xor X(329) xor X(331) xor X(332) xor X(333) xor X(334) xor X(335) xor X(337) xor X(338) xor X(339) xor X(341) xor X(342) xor X(345) xor X(346) xor X(350) xor X(351) xor X(352) xor X(353) xor X(356) xor X(360) xor X(363) xor X(364) xor X(366) xor X(367) xor X(368) xor X(376) xor X(377) xor X(380) xor X(384) xor X(385) xor X(387) xor X(388) xor X(392) xor X(393) xor X(394) xor X(395) xor X(396) xor X(400) xor X(401) xor X(406) xor X(407) xor X(410) xor X(411) xor X(413) xor X(415) xor X(417) xor X(418) xor X(419) xor X(421) xor X(424) xor X(427) xor X(430) xor X(432) xor X(439) xor X(441) xor X(442) xor X(443) xor X(446) xor X(447) xor X(448) xor X(449) xor X(451) xor X(453) xor X(454) xor X(459) xor X(460) xor X(461) xor X(462) xor X(464) xor X(465) xor X(467) xor X(469) xor X(472) xor X(473) xor X(474) xor X(475) xor X(476) xor X(480) xor X(486) xor X(487) xor X(493) xor X(494) xor X(496) xor X(499) xor X(503) xor X(505) xor X(508) xor X(509));
R_n(18) <= (R(0) xor R(6) xor R(7) xor R(9) xor R(12) xor R(16) xor R(18) xor R(21) xor R(22) xor X(1) xor X(3) xor X(4) xor X(5) xor X(6) xor X(7) xor X(8) xor X(9) xor X(10) xor X(11) xor X(12) xor X(13) xor X(14) xor X(17) xor X(20) xor X(21) xor X(23) xor X(24) xor X(25) xor X(28) xor X(35) xor X(37) xor X(38) xor X(39) xor X(40) xor X(42) xor X(44) xor X(45) xor X(46) xor X(49) xor X(50) xor X(51) xor X(52) xor X(55) xor X(56) xor X(57) xor X(60) xor X(61) xor X(63) xor X(64) xor X(65) xor X(66) xor X(67) xor X(68) xor X(70) xor X(75) xor X(78) xor X(79) xor X(82) xor X(83) xor X(86) xor X(87) xor X(88) xor X(89) xor X(91) xor X(92) xor X(93) xor X(97) xor X(100) xor X(101) xor X(102) xor X(104) xor X(105) xor X(107) xor X(110) xor X(111) xor X(112) xor X(113) xor X(115) xor X(118) xor X(121) xor X(122) xor X(123) xor X(126) xor X(127) xor X(128) xor X(132) xor X(136) xor X(137) xor X(138) xor X(140) xor X(142) xor X(144) xor X(151) xor X(152) xor X(154) xor X(155) xor X(156) xor X(158) xor X(164) xor X(169) xor X(171) xor X(172) xor X(173) xor X(174) xor X(175) xor X(176) xor X(177) xor X(182) xor X(183) xor X(186) xor X(188) xor X(190) xor X(192) xor X(196) xor X(197) xor X(199) xor X(200) xor X(201) xor X(202) xor X(203) xor X(204) xor X(205) xor X(210) xor X(211) xor X(213) xor X(214) xor X(215) xor X(217) xor X(219) xor X(220) xor X(224) xor X(225) xor X(226) xor X(230) xor X(231) xor X(232) xor X(234) xor X(235) xor X(239) xor X(241) xor X(242) xor X(243) xor X(245) xor X(246) xor X(247) xor X(250) xor X(253) xor X(255) xor X(256) xor X(258) xor X(259) xor X(261) xor X(264) xor X(267) xor X(268) xor X(269) xor X(270) xor X(272) xor X(277) xor X(278) xor X(280) xor X(281) xor X(285) xor X(289) xor X(292) xor X(296) xor X(298) xor X(301) xor X(302) xor X(303) xor X(304) xor X(305) xor X(307) xor X(313) xor X(314) xor X(315) xor X(318) xor X(319) xor X(320) xor X(326) xor X(327) xor X(328) xor X(329) xor X(330) xor X(332) xor X(333) xor X(334) xor X(335) xor X(336) xor X(338) xor X(339) xor X(340) xor X(342) xor X(343) xor X(346) xor X(347) xor X(351) xor X(352) xor X(353) xor X(354) xor X(357) xor X(361) xor X(364) xor X(365) xor X(367) xor X(368) xor X(369) xor X(377) xor X(378) xor X(381) xor X(385) xor X(386) xor X(388) xor X(389) xor X(393) xor X(394) xor X(395) xor X(396) xor X(397) xor X(401) xor X(402) xor X(407) xor X(408) xor X(411) xor X(412) xor X(414) xor X(416) xor X(418) xor X(419) xor X(420) xor X(422) xor X(425) xor X(428) xor X(431) xor X(433) xor X(440) xor X(442) xor X(443) xor X(444) xor X(447) xor X(448) xor X(449) xor X(450) xor X(452) xor X(454) xor X(455) xor X(460) xor X(461) xor X(462) xor X(463) xor X(465) xor X(466) xor X(468) xor X(470) xor X(473) xor X(474) xor X(475) xor X(476) xor X(477) xor X(481) xor X(487) xor X(488) xor X(494) xor X(495) xor X(497) xor X(500) xor X(504) xor X(506) xor X(509) xor X(510));
R_n(19) <= (R(0) xor R(1) xor R(7) xor R(8) xor R(10) xor R(13) xor R(17) xor R(19) xor R(22) xor R(23) xor X(2) xor X(4) xor X(5) xor X(6) xor X(7) xor X(8) xor X(9) xor X(10) xor X(11) xor X(12) xor X(13) xor X(14) xor X(15) xor X(18) xor X(21) xor X(22) xor X(24) xor X(25) xor X(26) xor X(29) xor X(36) xor X(38) xor X(39) xor X(40) xor X(41) xor X(43) xor X(45) xor X(46) xor X(47) xor X(50) xor X(51) xor X(52) xor X(53) xor X(56) xor X(57) xor X(58) xor X(61) xor X(62) xor X(64) xor X(65) xor X(66) xor X(67) xor X(68) xor X(69) xor X(71) xor X(76) xor X(79) xor X(80) xor X(83) xor X(84) xor X(87) xor X(88) xor X(89) xor X(90) xor X(92) xor X(93) xor X(94) xor X(98) xor X(101) xor X(102) xor X(103) xor X(105) xor X(106) xor X(108) xor X(111) xor X(112) xor X(113) xor X(114) xor X(116) xor X(119) xor X(122) xor X(123) xor X(124) xor X(127) xor X(128) xor X(129) xor X(133) xor X(137) xor X(138) xor X(139) xor X(141) xor X(143) xor X(145) xor X(152) xor X(153) xor X(155) xor X(156) xor X(157) xor X(159) xor X(165) xor X(170) xor X(172) xor X(173) xor X(174) xor X(175) xor X(176) xor X(177) xor X(178) xor X(183) xor X(184) xor X(187) xor X(189) xor X(191) xor X(193) xor X(197) xor X(198) xor X(200) xor X(201) xor X(202) xor X(203) xor X(204) xor X(205) xor X(206) xor X(211) xor X(212) xor X(214) xor X(215) xor X(216) xor X(218) xor X(220) xor X(221) xor X(225) xor X(226) xor X(227) xor X(231) xor X(232) xor X(233) xor X(235) xor X(236) xor X(240) xor X(242) xor X(243) xor X(244) xor X(246) xor X(247) xor X(248) xor X(251) xor X(254) xor X(256) xor X(257) xor X(259) xor X(260) xor X(262) xor X(265) xor X(268) xor X(269) xor X(270) xor X(271) xor X(273) xor X(278) xor X(279) xor X(281) xor X(282) xor X(286) xor X(290) xor X(293) xor X(297) xor X(299) xor X(302) xor X(303) xor X(304) xor X(305) xor X(306) xor X(308) xor X(314) xor X(315) xor X(316) xor X(319) xor X(320) xor X(321) xor X(327) xor X(328) xor X(329) xor X(330) xor X(331) xor X(333) xor X(334) xor X(335) xor X(336) xor X(337) xor X(339) xor X(340) xor X(341) xor X(343) xor X(344) xor X(347) xor X(348) xor X(352) xor X(353) xor X(354) xor X(355) xor X(358) xor X(362) xor X(365) xor X(366) xor X(368) xor X(369) xor X(370) xor X(378) xor X(379) xor X(382) xor X(386) xor X(387) xor X(389) xor X(390) xor X(394) xor X(395) xor X(396) xor X(397) xor X(398) xor X(402) xor X(403) xor X(408) xor X(409) xor X(412) xor X(413) xor X(415) xor X(417) xor X(419) xor X(420) xor X(421) xor X(423) xor X(426) xor X(429) xor X(432) xor X(434) xor X(441) xor X(443) xor X(444) xor X(445) xor X(448) xor X(449) xor X(450) xor X(451) xor X(453) xor X(455) xor X(456) xor X(461) xor X(462) xor X(463) xor X(464) xor X(466) xor X(467) xor X(469) xor X(471) xor X(474) xor X(475) xor X(476) xor X(477) xor X(478) xor X(482) xor X(488) xor X(489) xor X(495) xor X(496) xor X(498) xor X(501) xor X(505) xor X(507) xor X(510) xor X(511));
R_n(20) <= (R(0) xor R(1) xor R(2) xor R(4) xor R(5) xor R(6) xor R(7) xor R(8) xor R(9) xor R(12) xor R(13) xor R(15) xor R(19) xor R(20) xor R(21) xor R(22) xor X(0) xor X(4) xor X(5) xor X(9) xor X(12) xor X(13) xor X(15) xor X(19) xor X(22) xor X(25) xor X(26) xor X(27) xor X(29) xor X(31) xor X(32) xor X(34) xor X(36) xor X(38) xor X(40) xor X(42) xor X(44) xor X(47) xor X(49) xor X(51) xor X(54) xor X(56) xor X(57) xor X(60) xor X(64) xor X(68) xor X(72) xor X(73) xor X(81) xor X(83) xor X(84) xor X(86) xor X(87) xor X(88) xor X(90) xor X(93) xor X(94) xor X(95) xor X(97) xor X(98) xor X(100) xor X(102) xor X(106) xor X(109) xor X(112) xor X(114) xor X(115) xor X(117) xor X(118) xor X(119) xor X(120) xor X(125) xor X(126) xor X(127) xor X(128) xor X(129) xor X(130) xor X(131) xor X(132) xor X(133) xor X(134) xor X(137) xor X(139) xor X(142) xor X(144) xor X(148) xor X(149) xor X(151) xor X(155) xor X(161) xor X(163) xor X(164) xor X(165) xor X(171) xor X(173) xor X(174) xor X(176) xor X(178) xor X(179) xor X(182) xor X(183) xor X(184) xor X(187) xor X(188) xor X(191) xor X(193) xor X(196) xor X(198) xor X(200) xor X(201) xor X(202) xor X(206) xor X(208) xor X(211) xor X(213) xor X(214) xor X(215) xor X(216) xor X(217) xor X(218) xor X(220) xor X(221) xor X(222) xor X(223) xor X(224) xor X(225) xor X(226) xor X(227) xor X(228) xor X(229) xor X(230) xor X(231) xor X(232) xor X(233) xor X(234) xor X(235) xor X(240) xor X(241) xor X(246) xor X(251) xor X(254) xor X(255) xor X(259) xor X(262) xor X(263) xor X(264) xor X(265) xor X(269) xor X(270) xor X(271) xor X(272) xor X(273) xor X(275) xor X(278) xor X(280) xor X(281) xor X(282) xor X(283) xor X(285) xor X(286) xor X(288) xor X(292) xor X(295) xor X(296) xor X(297) xor X(300) xor X(303) xor X(305) xor X(306) xor X(307) xor X(310) xor X(311) xor X(312) xor X(313) xor X(315) xor X(316) xor X(319) xor X(320) xor X(321) xor X(323) xor X(324) xor X(326) xor X(333) xor X(337) xor X(339) xor X(340) xor X(341) xor X(343) xor X(345) xor X(346) xor X(348) xor X(349) xor X(350) xor X(352) xor X(353) xor X(358) xor X(361) xor X(363) xor X(364) xor X(365) xor X(366) xor X(367) xor X(372) xor X(373) xor X(374) xor X(375) xor X(380) xor X(382) xor X(383) xor X(384) xor X(385) xor X(386) xor X(387) xor X(388) xor X(392) xor X(393) xor X(394) xor X(396) xor X(397) xor X(398) xor X(399) xor X(400) xor X(401) xor X(402) xor X(403) xor X(404) xor X(406) xor X(407) xor X(408) xor X(410) xor X(413) xor X(416) xor X(418) xor X(421) xor X(423) xor X(424) xor X(426) xor X(428) xor X(429) xor X(430) xor X(431) xor X(436) xor X(438) xor X(439) xor X(440) xor X(441) xor X(442) xor X(444) xor X(450) xor X(451) xor X(456) xor X(462) xor X(463) xor X(464) xor X(465) xor X(466) xor X(470) xor X(471) xor X(472) xor X(477) xor X(482) xor X(483) xor X(485) xor X(486) xor X(487) xor X(488) xor X(489) xor X(490) xor X(492) xor X(493) xor X(494) xor X(495) xor X(496) xor X(497) xor X(500) xor X(501) xor X(503) xor X(507) xor X(508) xor X(509) xor X(510));
R_n(21) <= (R(1) xor R(2) xor R(3) xor R(4) xor R(8) xor R(9) xor R(10) xor R(11) xor R(12) xor R(15) xor R(16) xor R(18) xor R(19) xor R(20) xor X(0) xor X(1) xor X(3) xor X(4) xor X(5) xor X(7) xor X(8) xor X(11) xor X(13) xor X(20) xor X(26) xor X(27) xor X(28) xor X(29) xor X(31) xor X(33) xor X(34) xor X(35) xor X(36) xor X(38) xor X(43) xor X(45) xor X(46) xor X(49) xor X(50) xor X(53) xor X(55) xor X(56) xor X(57) xor X(59) xor X(60) xor X(61) xor X(62) xor X(63) xor X(64) xor X(66) xor X(67) xor X(70) xor X(74) xor X(77) xor X(80) xor X(82) xor X(83) xor X(84) xor X(86) xor X(88) xor X(94) xor X(95) xor X(96) xor X(97) xor X(100) xor X(101) xor X(104) xor X(110) xor X(115) xor X(116) xor X(120) xor X(121) xor X(123) xor X(124) xor X(128) xor X(129) xor X(130) xor X(134) xor X(135) xor X(137) xor X(143) xor X(145) xor X(146) xor X(148) xor X(150) xor X(151) xor X(152) xor X(153) xor X(154) xor X(155) xor X(157) xor X(158) xor X(160) xor X(161) xor X(162) xor X(163) xor X(172) xor X(174) xor X(179) xor X(180) xor X(182) xor X(184) xor X(187) xor X(188) xor X(189) xor X(190) xor X(191) xor X(193) xor X(196) xor X(197) xor X(200) xor X(201) xor X(202) xor X(204) xor X(205) xor X(208) xor X(209) xor X(211) xor X(215) xor X(216) xor X(217) xor X(220) xor X(221) xor X(222) xor X(226) xor X(227) xor X(228) xor X(232) xor X(233) xor X(234) xor X(237) xor X(240) xor X(241) xor X(242) xor X(243) xor X(244) xor X(245) xor X(246) xor X(248) xor X(249) xor X(251) xor X(254) xor X(255) xor X(256) xor X(257) xor X(258) xor X(259) xor X(261) xor X(262) xor X(263) xor X(270) xor X(271) xor X(272) xor X(275) xor X(276) xor X(278) xor X(282) xor X(283) xor X(284) xor X(285) xor X(288) xor X(289) xor X(291) xor X(292) xor X(293) xor X(294) xor X(295) xor X(301) xor X(306) xor X(307) xor X(308) xor X(309) xor X(310) xor X(314) xor X(316) xor X(319) xor X(320) xor X(321) xor X(323) xor X(325) xor X(326) xor X(327) xor X(328) xor X(329) xor X(330) xor X(331) xor X(332) xor X(333) xor X(335) xor X(336) xor X(339) xor X(340) xor X(341) xor X(343) xor X(347) xor X(349) xor X(351) xor X(352) xor X(353) xor X(355) xor X(356) xor X(358) xor X(361) xor X(362) xor X(366) xor X(367) xor X(368) xor X(369) xor X(370) xor X(371) xor X(372) xor X(376) xor X(379) xor X(381) xor X(382) xor X(383) xor X(387) xor X(388) xor X(389) xor X(390) xor X(391) xor X(392) xor X(397) xor X(398) xor X(399) xor X(403) xor X(404) xor X(405) xor X(406) xor X(411) xor X(417) xor X(419) xor X(420) xor X(423) xor X(424) xor X(425) xor X(426) xor X(428) xor X(430) xor X(432) xor X(433) xor X(435) xor X(436) xor X(437) xor X(438) xor X(442) xor X(443) xor X(446) xor X(449) xor X(451) xor X(454) xor X(463) xor X(464) xor X(465) xor X(468) xor X(472) xor X(473) xor X(475) xor X(476) xor X(479) xor X(482) xor X(483) xor X(484) xor X(485) xor X(489) xor X(490) xor X(491) xor X(492) xor X(496) xor X(497) xor X(498) xor X(499) xor X(500) xor X(503) xor X(504) xor X(506) xor X(507) xor X(508));
R_n(22) <= (R(2) xor R(3) xor R(4) xor R(5) xor R(9) xor R(10) xor R(11) xor R(12) xor R(13) xor R(16) xor R(17) xor R(19) xor R(20) xor R(21) xor X(1) xor X(2) xor X(4) xor X(5) xor X(6) xor X(8) xor X(9) xor X(12) xor X(14) xor X(21) xor X(27) xor X(28) xor X(29) xor X(30) xor X(32) xor X(34) xor X(35) xor X(36) xor X(37) xor X(39) xor X(44) xor X(46) xor X(47) xor X(50) xor X(51) xor X(54) xor X(56) xor X(57) xor X(58) xor X(60) xor X(61) xor X(62) xor X(63) xor X(64) xor X(65) xor X(67) xor X(68) xor X(71) xor X(75) xor X(78) xor X(81) xor X(83) xor X(84) xor X(85) xor X(87) xor X(89) xor X(95) xor X(96) xor X(97) xor X(98) xor X(101) xor X(102) xor X(105) xor X(111) xor X(116) xor X(117) xor X(121) xor X(122) xor X(124) xor X(125) xor X(129) xor X(130) xor X(131) xor X(135) xor X(136) xor X(138) xor X(144) xor X(146) xor X(147) xor X(149) xor X(151) xor X(152) xor X(153) xor X(154) xor X(155) xor X(156) xor X(158) xor X(159) xor X(161) xor X(162) xor X(163) xor X(164) xor X(173) xor X(175) xor X(180) xor X(181) xor X(183) xor X(185) xor X(188) xor X(189) xor X(190) xor X(191) xor X(192) xor X(194) xor X(197) xor X(198) xor X(201) xor X(202) xor X(203) xor X(205) xor X(206) xor X(209) xor X(210) xor X(212) xor X(216) xor X(217) xor X(218) xor X(221) xor X(222) xor X(223) xor X(227) xor X(228) xor X(229) xor X(233) xor X(234) xor X(235) xor X(238) xor X(241) xor X(242) xor X(243) xor X(244) xor X(245) xor X(246) xor X(247) xor X(249) xor X(250) xor X(252) xor X(255) xor X(256) xor X(257) xor X(258) xor X(259) xor X(260) xor X(262) xor X(263) xor X(264) xor X(271) xor X(272) xor X(273) xor X(276) xor X(277) xor X(279) xor X(283) xor X(284) xor X(285) xor X(286) xor X(289) xor X(290) xor X(292) xor X(293) xor X(294) xor X(295) xor X(296) xor X(302) xor X(307) xor X(308) xor X(309) xor X(310) xor X(311) xor X(315) xor X(317) xor X(320) xor X(321) xor X(322) xor X(324) xor X(326) xor X(327) xor X(328) xor X(329) xor X(330) xor X(331) xor X(332) xor X(333) xor X(334) xor X(336) xor X(337) xor X(340) xor X(341) xor X(342) xor X(344) xor X(348) xor X(350) xor X(352) xor X(353) xor X(354) xor X(356) xor X(357) xor X(359) xor X(362) xor X(363) xor X(367) xor X(368) xor X(369) xor X(370) xor X(371) xor X(372) xor X(373) xor X(377) xor X(380) xor X(382) xor X(383) xor X(384) xor X(388) xor X(389) xor X(390) xor X(391) xor X(392) xor X(393) xor X(398) xor X(399) xor X(400) xor X(404) xor X(405) xor X(406) xor X(407) xor X(412) xor X(418) xor X(420) xor X(421) xor X(424) xor X(425) xor X(426) xor X(427) xor X(429) xor X(431) xor X(433) xor X(434) xor X(436) xor X(437) xor X(438) xor X(439) xor X(443) xor X(444) xor X(447) xor X(450) xor X(452) xor X(455) xor X(464) xor X(465) xor X(466) xor X(469) xor X(473) xor X(474) xor X(476) xor X(477) xor X(480) xor X(483) xor X(484) xor X(485) xor X(486) xor X(490) xor X(491) xor X(492) xor X(493) xor X(497) xor X(498) xor X(499) xor X(500) xor X(501) xor X(504) xor X(505) xor X(507) xor X(508) xor X(509));
R_n(23) <= (R(3) xor R(4) xor R(5) xor R(6) xor R(10) xor R(11) xor R(12) xor R(13) xor R(14) xor R(17) xor R(18) xor R(20) xor R(21) xor R(22) xor X(2) xor X(3) xor X(5) xor X(6) xor X(7) xor X(9) xor X(10) xor X(13) xor X(15) xor X(22) xor X(28) xor X(29) xor X(30) xor X(31) xor X(33) xor X(35) xor X(36) xor X(37) xor X(38) xor X(40) xor X(45) xor X(47) xor X(48) xor X(51) xor X(52) xor X(55) xor X(57) xor X(58) xor X(59) xor X(61) xor X(62) xor X(63) xor X(64) xor X(65) xor X(66) xor X(68) xor X(69) xor X(72) xor X(76) xor X(79) xor X(82) xor X(84) xor X(85) xor X(86) xor X(88) xor X(90) xor X(96) xor X(97) xor X(98) xor X(99) xor X(102) xor X(103) xor X(106) xor X(112) xor X(117) xor X(118) xor X(122) xor X(123) xor X(125) xor X(126) xor X(130) xor X(131) xor X(132) xor X(136) xor X(137) xor X(139) xor X(145) xor X(147) xor X(148) xor X(150) xor X(152) xor X(153) xor X(154) xor X(155) xor X(156) xor X(157) xor X(159) xor X(160) xor X(162) xor X(163) xor X(164) xor X(165) xor X(174) xor X(176) xor X(181) xor X(182) xor X(184) xor X(186) xor X(189) xor X(190) xor X(191) xor X(192) xor X(193) xor X(195) xor X(198) xor X(199) xor X(202) xor X(203) xor X(204) xor X(206) xor X(207) xor X(210) xor X(211) xor X(213) xor X(217) xor X(218) xor X(219) xor X(222) xor X(223) xor X(224) xor X(228) xor X(229) xor X(230) xor X(234) xor X(235) xor X(236) xor X(239) xor X(242) xor X(243) xor X(244) xor X(245) xor X(246) xor X(247) xor X(248) xor X(250) xor X(251) xor X(253) xor X(256) xor X(257) xor X(258) xor X(259) xor X(260) xor X(261) xor X(263) xor X(264) xor X(265) xor X(272) xor X(273) xor X(274) xor X(277) xor X(278) xor X(280) xor X(284) xor X(285) xor X(286) xor X(287) xor X(290) xor X(291) xor X(293) xor X(294) xor X(295) xor X(296) xor X(297) xor X(303) xor X(308) xor X(309) xor X(310) xor X(311) xor X(312) xor X(316) xor X(318) xor X(321) xor X(322) xor X(323) xor X(325) xor X(327) xor X(328) xor X(329) xor X(330) xor X(331) xor X(332) xor X(333) xor X(334) xor X(335) xor X(337) xor X(338) xor X(341) xor X(342) xor X(343) xor X(345) xor X(349) xor X(351) xor X(353) xor X(354) xor X(355) xor X(357) xor X(358) xor X(360) xor X(363) xor X(364) xor X(368) xor X(369) xor X(370) xor X(371) xor X(372) xor X(373) xor X(374) xor X(378) xor X(381) xor X(383) xor X(384) xor X(385) xor X(389) xor X(390) xor X(391) xor X(392) xor X(393) xor X(394) xor X(399) xor X(400) xor X(401) xor X(405) xor X(406) xor X(407) xor X(408) xor X(413) xor X(419) xor X(421) xor X(422) xor X(425) xor X(426) xor X(427) xor X(428) xor X(430) xor X(432) xor X(434) xor X(435) xor X(437) xor X(438) xor X(439) xor X(440) xor X(444) xor X(445) xor X(448) xor X(451) xor X(453) xor X(456) xor X(465) xor X(466) xor X(467) xor X(470) xor X(474) xor X(475) xor X(477) xor X(478) xor X(481) xor X(484) xor X(485) xor X(486) xor X(487) xor X(491) xor X(492) xor X(493) xor X(494) xor X(498) xor X(499) xor X(500) xor X(501) xor X(502) xor X(505) xor X(506) xor X(508) xor X(509) xor X(510));

end functional;
