// import lynxTypes::*;

// Replace the Streaming Inputs with simple bit inputs for easier testing 

module icrc(
    // Networking interface - Incoming and outgoing traffic - for ease of use, revert back to simple bitfields 
    AXI4S.s m_axis_rx, 
    AXI4S.m m_axis_tx, 

    // Incoming clock and reset
    input logic nclk, 
    input logic nresetn
);


//////////////////////////////////////////////////////////////////////////////////////
//
// Definition of data types 
//
//////////////////////////////////////////////////////////////////////////////////////

// 512 Bit Data Type to hold the incoming words 
typedef logic [511:0] DataWord;

// 64 Bit Data Type to hold the incoming keep value
typedef logic [63:0] KeepWord; 

// 16 Bit Data Type to determine which of the CRC32 pipeline-stages need to be used 
typedef logic [15:0] CRC32ValidStages; 

// 32 Bit Data Type to hold the CRC values
typedef logic [31:0] CRCWord; 

// SubKeepWord for Probing only 
typedef logic [3:0] SubKeepWord; 

// CounterWord for CRC32 stages
typedef logic [3:0] CRC32CounterWord;  


///////////////////////////////////////////////////////////////////////////////////////
// 
// Definition of registers for the Pipeline Stages
//
///////////////////////////////////////////////////////////////////////////////////////

// Regs for the masking stage 
logic stage_masking_valid; 
DataWord stage_masking_data; 
DataWord stage_masking_masked_data; 
KeepWord stage_masking_keep; 
logic stage_masking_last; 
logic stage_crc_follow_up_word; 
CRCWord stage_masking_crc_seed; 

// Regs for the CRC32-pipeline stages 
logic stage_crc32_valid[16]; 
DataWord stage_crc32_data_bypass[16]; 
DataWord stage_crc32_masked_data[16]; 
CRCWord stage_crc32_crc[16]; 
KeepWord stage_crc32_keep[16];
logic stage_crc32_last[16]; 
CRC32ValidStages stage_crc32_valid_stages[16];  
SubKeepWord stage_crc32_keep_stage[16]; 
logic stage_crc32_early_done; 
CRC32CounterWord stage_crc32_counter_word; 


// Regs for the CRC512-pipeline stage 
logic stage_crc512_valid;
DataWord stage_crc512_data_bypass; 
DataWord stage_crc512_masked_data; 
CRCWord stage_crc512_crc; 
KeepWord stage_crc512_keep; 
logic stage_crc512_last; 

// Regs for the CRC320-pipeline stage 
logic stage_crc320_valid; 
DataWord stage_crc320_data_bypass; 
DataWord stage_crc320_masked_data; 
CRCWord stage_crc320_crc; 
KeepWord stage_crc320_keep; 
logic stage_crc320_last; 

// Regs for the pipeline-join-stage 
logic stage_join_valid; 
DataWord stage_join_data; 
CRCWord stage_join_crc; 
KeepWord stage_join_keep; 
logic stage_join_last; 

// Regs for the reinsertion stage 
logic stage_reinsertion_valid; 
DataWord stage_reinsertion_data; 
CRCWord stage_reinsertion_crc; 
KeepWord stage_reinsertion_keep; 
logic stage_reinsertion_last; 

// Regs for the last add-word stage 
logic stage_add_word_valid; 
DataWord stage_add_word_data;
CRCWord stage_add_word_crc; 
KeepWord stage_add_word_keep;
logic stage_add_word_last; 

// Wires from the pipeline to the final buffer-FIFO 
DataWord pipeline_to_fifo_data; 
KeepWord pipeline_to_fifo_keep; 
logic pipeline_to_fifo_last; 
logic pipeline_to_fifo_valid; 
logic pipeline_to_fifo_reset; 
logic empty_output; 

// Register for stalling the pipeline 
logic stall_pipeline; 

// Register for controlling the output 
logic switch_output; 

// Bitmask for masking away the the unrequired fields of the incoming data 
DataWord bitmask; 

// Signal for assigning the ready signal at output 
logic halffull_signal; 
logic full_signal; 

// Define alias for CRC-seed and CRC-input data for CRC512 to avoid long lines that break the editor 
DataWord d; 
CRCWord c; 

// Test Probe to see if the CRC32 pipeline after [0] is activated at all 
logic crc32_test_probe; 
CRCWord crc32_data_probe[16]; 
CRCWord crc32_seed_probe[16]; 
logic crc32_in_flight; 
logic crc32_in_flight_comb; 

// Assign the initial CRC-inputs
assign d = stage_crc_follow_up_word ? stage_masking_data : stage_masking_masked_data; 
assign c = stage_crc_follow_up_word ? stage_crc512_crc : 32'hdebb20e3; 

// Assign the crc32-stage keeps 
assign stage_crc32_keep_stage[0] = stage_masking_keep[3:0]; 
assign stage_crc32_keep_stage[1] = stage_crc32_keep[0][7:4]; 
assign stage_crc32_keep_stage[2] = stage_crc32_keep[1][11:8]; 
assign stage_crc32_keep_stage[3] = stage_crc32_keep[2][15:12]; 
assign stage_crc32_keep_stage[4] = stage_crc32_keep[3][19:16]; 
assign stage_crc32_keep_stage[5] = stage_crc32_keep[4][23:20]; 
assign stage_crc32_keep_stage[6] = stage_crc32_keep[5][27:24]; 
assign stage_crc32_keep_stage[7] = stage_crc32_keep[6][31:28];
assign stage_crc32_keep_stage[8] = stage_crc32_keep[7][35:32];
assign stage_crc32_keep_stage[9] = stage_crc32_keep[8][39:36]; 
assign stage_crc32_keep_stage[10] = stage_crc32_keep[9][43:40]; 
assign stage_crc32_keep_stage[11] = stage_crc32_keep[10][47:44];
assign stage_crc32_keep_stage[12] = stage_crc32_keep[11][51:48]; 
assign stage_crc32_keep_stage[13] = stage_crc32_keep[12][55:52];
assign stage_crc32_keep_stage[14] = stage_crc32_keep[13][59:56]; 
assign stage_crc32_keep_stage[15] = stage_crc32_keep[14][63:60];

// Assign the calculation of the crc32_in_flight_comb signal that goes high in the very clock cycle when a CRC32-candidate is detected 
assign crc32_in_flight_comb = crc32_in_flight || ((stage_masking_keep != 64'hffffffffffffffff) && (stage_masking_keep != 64'h000000ffffffffff) && (stage_masking_keep != 64'h0));



/////////////////////////////////////////////////////////////////////////////////////////////
//
// Assignment of d for CRC-calculation to stage_1_bitmasked data
//
/////////////////////////////////////////////////////////////////////////////////////////////

always_ff @(posedge nclk) begin

    // Reset of all stage signals 
    if(!nresetn) begin 
        // Reset of the masking stage 
        stage_masking_valid <= 1'b0; 
        stage_masking_data <= 512'b0;
        stage_masking_masked_data <= 512'b0; 
        stage_masking_keep <= 64'b0; 
        stage_masking_last <= 1'b0; 
        stage_crc_follow_up_word <= 1'b0; 
        stage_masking_crc_seed <= 32'b0; 

        // Reset of the CRC32-pipeline stages in parallel 
        for(integer pipeline_stage = 0; pipeline_stage < 16; pipeline_stage++) begin
            stage_crc32_valid[pipeline_stage] <= 1'b0; 
            stage_crc32_data_bypass[pipeline_stage] <= 512'b0; 
            stage_crc32_masked_data[pipeline_stage] <= 512'b0;
            stage_crc32_crc[pipeline_stage] <= 32'b0;
            stage_crc32_keep[pipeline_stage] <= 64'b0;
            stage_crc32_last[pipeline_stage] <= 1'b0; 
            stage_crc32_valid_stages[pipeline_stage] <= 32'b0;
            crc32_data_probe[pipeline_stage] <= 32'b0; 
            crc32_seed_probe[pipeline_stage] <= 32'b0;  
        end

        stage_crc32_counter_word <= 4'b0; 
        stage_crc32_early_done <= 1'b0; 

        // Reset of the CRC512-pipeline stage
        stage_crc512_valid <= 1'b0; 
        stage_crc512_data_bypass <= 512'b0;
        stage_crc512_masked_data <= 512'b0; 
        stage_crc512_crc <= 32'b0;
        stage_crc512_keep <= 64'b0; 
        stage_crc512_last <= 1'b0; 

        // Reset of the CRC320-pipeline stage 
        stage_crc320_valid <= 1'b0; 
        stage_crc320_data_bypass <= 512'b0; 
        stage_crc320_masked_data <= 512'b0; 
        stage_crc320_crc <= 32'b0;
        stage_crc320_keep <= 64'b0; 
        stage_crc320_last <= 1'b0; 

        // Reset of the join pipeline stage 
        stage_join_valid <= 1'b0; 
        stage_join_data <= 512'b0; 
        stage_join_crc <= 32'b0; 
        stage_join_keep <= 64'b0; 
        stage_join_last <= 1'b0; 

        // Reset of the reinsertion pipeline stage 
        stage_reinsertion_valid <= 1'b0; 
        stage_reinsertion_data <= 512'b0; 
        stage_reinsertion_crc <= 32'b0; 
        stage_reinsertion_keep <= 64'b0; 
        stage_reinsertion_last <= 1'b0;  

        // Reset of the Add-Word-Stage 
        stage_add_word_valid <= 1'b0; 
        stage_add_word_data <= 512'b0; 
        stage_add_word_crc <= 32'b0; 
        stage_add_word_keep <= 64'b0; 
        stage_add_word_last <= 1'b0; 

        // Reset of the register for stalling the pipeline 
        stall_pipeline <= 1'b0; 
        crc32_in_flight <= 1'b0; 

        // Reset of the register for switching the output 
        switch_output <= 1'b0; 

        // Set-Up of the bitmask 
        bitmask[351:0] <= 352'h0000000000000000000000ff00000000ffff0000000000000000000000000000ffff00ff000000000000ff00; 
        bitmask[511:352] <= 160'b0; 

        // Reset the test probe 
        crc32_test_probe <= 1'b0; 

    end else begin

        /////////////////////////////////////////////////////////////////////
        //
        // STAGE 1: LOADING AND BITMASKING
        //
        /////////////////////////////////////////////////////////////////////
        
        if(~halffull_signal & ~crc32_in_flight_comb & ~full_signal) begin 
            // Forward direct signals: valid, last, keep, data 
            stage_masking_valid <= m_axis_rx.tvalid;
            stage_masking_last <= m_axis_rx.tlast;
            stage_masking_keep <= m_axis_rx.tkeep;
            stage_masking_data <= m_axis_rx.tdata;

            // If input is valid, load and mask data - else it's just 0s 
            if(m_axis_rx.tvalid) begin 
                // Only mask the first word (only one with Header Fields)
                if(stage_crc_follow_up_word == 0) begin 
                    stage_masking_masked_data <= m_axis_rx.tdata | bitmask; 

                    // Set the initial crc-value to debb20e3 (CRC of the imaginary leading GRH) and insert to the correct CRC-pipeline 
                    stage_masking_crc_seed <= 32'hdebb20e3; 

                    // if(m_axis_rx.tkeep == 64'hffffffffffffffff) begin 
                    //     // Full 512-bit word, can go to CRC512 pipeline
                    //     stage_crc512_crc <= 32'hdebb20e3; 
                    // end else if(m_axis_rx.tkeep == 64'h000000ffffffffff) begin 
                    //     // 320-bit word, can go to CRC320 pipeline 
                    //     stage_crc320_crc <= 32'hdebb20e3; 
                    // end else begin 
                    //     // Other 4-byte aligned word, must go to CRC32 pipeline 
                    //     stage_crc32_crc <= 32'hdebb20e3; 
                    // end 
                end else begin
                    stage_masking_masked_data <= m_axis_rx.tdata; 
                    
                    // Use the crc512 output, since in many-word cases all except the last one will be 512 bit anyways
                    stage_masking_crc_seed <= stage_crc512_crc; 
                end 
            end
        end else begin 
            // If the pipeline is full, stall the input
            stage_masking_valid <= 1'b0;
            stage_masking_keep <= 64'b0;
            stage_masking_data <= 512'b0;
            stage_masking_last <= 1'b0;
        end 


        ///////////////////////////////////////////////////////////////////////
        //
        // STAGE 2: CRC-Calculation 
        //
        ///////////////////////////////////////////////////////////////////////

        // Depending on the incoming keep-value, choose on of the three available CRC-pipelines (512, 320 or 32 Bits)
        if(stage_masking_valid) begin 

            // Calculate the word indicator
            if(!stage_masking_last) begin
                stage_crc_follow_up_word <= 1; 
                // stage_crc32_masked_data[0] <= stage_masking_data;  
            end else begin 
                stage_crc_follow_up_word <= 0;
                // stage_crc32_masked_data[0] <= stage_masking_masked_data; 
            end

            if(stage_masking_keep == 64'hffffffffffffffff) begin

                // === CRC512 ===

                // Forward direct signals: valid, last, keep, data_bypass
                stage_crc512_valid <= stage_masking_valid; 
                stage_crc512_last <= stage_masking_last; 
                stage_crc512_keep <= stage_masking_keep;
                stage_crc512_data_bypass <= stage_masking_data; 

                // Reset all other signals of the parallel CRC pipelines 
                stage_crc320_valid <= 1'b0;
                stage_crc320_last <= 1'b0; 
                stage_crc320_keep <= 64'b0; 
                stage_crc320_data_bypass <= 512'b0; 
                stage_crc320_crc <= 32'b0; 

                for(integer pipeline_stage = 0; pipeline_stage < 16; pipeline_stage++) begin
                    stage_crc32_valid[pipeline_stage] <= 1'b0; 
                    stage_crc32_last[pipeline_stage] <= 1'b0; 
                    stage_crc32_keep[pipeline_stage] <= 64'b0; 
                    stage_crc32_data_bypass[pipeline_stage] <= 512'b0; 
                    stage_crc32_crc[pipeline_stage] <= 32'b0; 
                end  


                // Bitwise calculation of the CRC512-value based on the bitmasked data and the CRC-seed. 
                stage_crc512_crc[31] <= d[511-511] ^ d[511-510] ^ d[511-508] ^ d[511-507] ^ d[511-506] ^ d[511-502] ^ d[511-501] ^ d[511-500] ^ d[511-495] ^ d[511-494] ^ d[511-493] ^ d[511-492] ^ d[511-491] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-486] ^ d[511-483] ^ d[511-482] ^ d[511-481] ^ d[511-480] ^ d[511-479] ^ d[511-477] ^ d[511-476] ^ d[511-472] ^ d[511-470] ^ d[511-468] ^ d[511-465] ^ d[511-464] ^ d[511-462] ^ d[511-461] ^ d[511-458] ^ d[511-452] ^ d[511-450] ^ d[511-449] ^ d[511-448] ^ d[511-444] ^ d[511-437] ^ d[511-436] ^ d[511-434] ^ d[511-433] ^ d[511-424] ^ d[511-422] ^ d[511-419] ^ d[511-418] ^ d[511-416] ^ d[511-414] ^ d[511-412] ^ d[511-409] ^ d[511-408] ^ d[511-407] ^ d[511-405] ^ d[511-404] ^ d[511-400] ^ d[511-399] ^ d[511-398] ^ d[511-396] ^ d[511-393] ^ d[511-392] ^ d[511-391] ^ d[511-390] ^ d[511-388] ^ d[511-387] ^ d[511-386] ^ d[511-381] ^ d[511-378] ^ d[511-376] ^ d[511-374] ^ d[511-372] ^ d[511-369] ^ d[511-368] ^ d[511-366] ^ d[511-363] ^ d[511-362] ^ d[511-359] ^ d[511-358] ^ d[511-357] ^ d[511-353] ^ d[511-349] ^ d[511-348] ^ d[511-347] ^ d[511-345] ^ d[511-344] ^ d[511-342] ^ d[511-341] ^ d[511-339] ^ d[511-338] ^ d[511-337] ^ d[511-335] ^ d[511-334] ^ d[511-333] ^ d[511-328] ^ d[511-327] ^ d[511-322] ^ d[511-321] ^ d[511-320] ^ d[511-319] ^ d[511-318] ^ d[511-317] ^ d[511-315] ^ d[511-312] ^ d[511-310] ^ d[511-309] ^ d[511-305] ^ d[511-303] ^ d[511-302] ^ d[511-300] ^ d[511-299] ^ d[511-298] ^ d[511-297] ^ d[511-296] ^ d[511-295] ^ d[511-294] ^ d[511-292] ^ d[511-290] ^ d[511-288] ^ d[511-287] ^ d[511-286] ^ d[511-283] ^ d[511-279] ^ d[511-277] ^ d[511-276] ^ d[511-274] ^ d[511-273] ^ d[511-269] ^ d[511-268] ^ d[511-265] ^ d[511-264] ^ d[511-261] ^ d[511-259] ^ d[511-257] ^ d[511-255] ^ d[511-252] ^ d[511-248] ^ d[511-243] ^ d[511-237] ^ d[511-234] ^ d[511-230] ^ d[511-228] ^ d[511-227] ^ d[511-226] ^ d[511-224] ^ d[511-216] ^ d[511-214] ^ d[511-212] ^ d[511-210] ^ d[511-209] ^ d[511-208] ^ d[511-207] ^ d[511-203] ^ d[511-202] ^ d[511-201] ^ d[511-199] ^ d[511-198] ^ d[511-197] ^ d[511-194] ^ d[511-193] ^ d[511-192] ^ d[511-191] ^ d[511-190] ^ d[511-188] ^ d[511-186] ^ d[511-183] ^ d[511-182] ^ d[511-172] ^ d[511-171] ^ d[511-170] ^ d[511-169] ^ d[511-167] ^ d[511-166] ^ d[511-162] ^ d[511-161] ^ d[511-158] ^ d[511-156] ^ d[511-155] ^ d[511-151] ^ d[511-149] ^ d[511-144] ^ d[511-143] ^ d[511-137] ^ d[511-136] ^ d[511-135] ^ d[511-134] ^ d[511-132] ^ d[511-128] ^ d[511-127] ^ d[511-126] ^ d[511-125] ^ d[511-123] ^ d[511-119] ^ d[511-118] ^ d[511-117] ^ d[511-116] ^ d[511-114] ^ d[511-113] ^ d[511-111] ^ d[511-110] ^ d[511-106] ^ d[511-104] ^ d[511-103] ^ d[511-101] ^ d[511-99] ^ d[511-98] ^ d[511-97] ^ d[511-96] ^ d[511-95] ^ d[511-94] ^ d[511-87] ^ d[511-85] ^ d[511-84] ^ d[511-83] ^ d[511-82] ^ d[511-81] ^ d[511-79] ^ d[511-73] ^ d[511-72] ^ d[511-68] ^ d[511-67] ^ d[511-66] ^ d[511-65] ^ d[511-63] ^ d[511-61] ^ d[511-60] ^ d[511-58] ^ d[511-55] ^ d[511-54] ^ d[511-53] ^ d[511-50] ^ d[511-48] ^ d[511-47] ^ d[511-45] ^ d[511-44] ^ d[511-37] ^ d[511-34] ^ d[511-32] ^ d[511-31] ^ d[511-30] ^ d[511-29] ^ d[511-28] ^ d[511-26] ^ d[511-25] ^ d[511-24] ^ d[511-16] ^ d[511-12] ^ d[511-10] ^ d[511-9] ^ d[511-6] ^ d[511-0] ^ c[31-0] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-6] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-20] ^ c[31-21] ^ c[31-22] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-30] ^ c[31-31];
                stage_crc512_crc[30] <= d[511-510] ^ d[511-509] ^ d[511-506] ^ d[511-503] ^ d[511-500] ^ d[511-496] ^ d[511-488] ^ d[511-487] ^ d[511-486] ^ d[511-484] ^ d[511-479] ^ d[511-478] ^ d[511-476] ^ d[511-473] ^ d[511-472] ^ d[511-471] ^ d[511-470] ^ d[511-469] ^ d[511-468] ^ d[511-466] ^ d[511-464] ^ d[511-463] ^ d[511-461] ^ d[511-459] ^ d[511-458] ^ d[511-453] ^ d[511-452] ^ d[511-451] ^ d[511-448] ^ d[511-445] ^ d[511-444] ^ d[511-438] ^ d[511-436] ^ d[511-435] ^ d[511-433] ^ d[511-425] ^ d[511-424] ^ d[511-423] ^ d[511-422] ^ d[511-420] ^ d[511-418] ^ d[511-417] ^ d[511-416] ^ d[511-415] ^ d[511-414] ^ d[511-413] ^ d[511-412] ^ d[511-410] ^ d[511-407] ^ d[511-406] ^ d[511-404] ^ d[511-401] ^ d[511-398] ^ d[511-397] ^ d[511-396] ^ d[511-394] ^ d[511-390] ^ d[511-389] ^ d[511-386] ^ d[511-382] ^ d[511-381] ^ d[511-379] ^ d[511-378] ^ d[511-377] ^ d[511-376] ^ d[511-375] ^ d[511-374] ^ d[511-373] ^ d[511-372] ^ d[511-370] ^ d[511-368] ^ d[511-367] ^ d[511-366] ^ d[511-364] ^ d[511-362] ^ d[511-360] ^ d[511-357] ^ d[511-354] ^ d[511-353] ^ d[511-350] ^ d[511-347] ^ d[511-346] ^ d[511-344] ^ d[511-343] ^ d[511-341] ^ d[511-340] ^ d[511-337] ^ d[511-336] ^ d[511-333] ^ d[511-329] ^ d[511-327] ^ d[511-323] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-313] ^ d[511-312] ^ d[511-311] ^ d[511-309] ^ d[511-306] ^ d[511-305] ^ d[511-304] ^ d[511-302] ^ d[511-301] ^ d[511-294] ^ d[511-293] ^ d[511-292] ^ d[511-291] ^ d[511-290] ^ d[511-289] ^ d[511-286] ^ d[511-284] ^ d[511-283] ^ d[511-280] ^ d[511-279] ^ d[511-278] ^ d[511-276] ^ d[511-275] ^ d[511-273] ^ d[511-270] ^ d[511-268] ^ d[511-266] ^ d[511-264] ^ d[511-262] ^ d[511-261] ^ d[511-260] ^ d[511-259] ^ d[511-258] ^ d[511-257] ^ d[511-256] ^ d[511-255] ^ d[511-253] ^ d[511-252] ^ d[511-249] ^ d[511-248] ^ d[511-244] ^ d[511-243] ^ d[511-238] ^ d[511-237] ^ d[511-235] ^ d[511-234] ^ d[511-231] ^ d[511-230] ^ d[511-229] ^ d[511-226] ^ d[511-225] ^ d[511-224] ^ d[511-217] ^ d[511-216] ^ d[511-215] ^ d[511-214] ^ d[511-213] ^ d[511-212] ^ d[511-211] ^ d[511-207] ^ d[511-204] ^ d[511-201] ^ d[511-200] ^ d[511-197] ^ d[511-195] ^ d[511-190] ^ d[511-189] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-184] ^ d[511-182] ^ d[511-173] ^ d[511-169] ^ d[511-168] ^ d[511-166] ^ d[511-163] ^ d[511-161] ^ d[511-159] ^ d[511-158] ^ d[511-157] ^ d[511-155] ^ d[511-152] ^ d[511-151] ^ d[511-150] ^ d[511-149] ^ d[511-145] ^ d[511-143] ^ d[511-138] ^ d[511-134] ^ d[511-133] ^ d[511-132] ^ d[511-129] ^ d[511-125] ^ d[511-124] ^ d[511-123] ^ d[511-120] ^ d[511-116] ^ d[511-115] ^ d[511-113] ^ d[511-112] ^ d[511-110] ^ d[511-107] ^ d[511-106] ^ d[511-105] ^ d[511-103] ^ d[511-102] ^ d[511-101] ^ d[511-100] ^ d[511-94] ^ d[511-88] ^ d[511-87] ^ d[511-86] ^ d[511-81] ^ d[511-80] ^ d[511-79] ^ d[511-74] ^ d[511-72] ^ d[511-69] ^ d[511-65] ^ d[511-64] ^ d[511-63] ^ d[511-62] ^ d[511-60] ^ d[511-59] ^ d[511-58] ^ d[511-56] ^ d[511-53] ^ d[511-51] ^ d[511-50] ^ d[511-49] ^ d[511-47] ^ d[511-46] ^ d[511-44] ^ d[511-38] ^ d[511-37] ^ d[511-35] ^ d[511-34] ^ d[511-33] ^ d[511-28] ^ d[511-27] ^ d[511-24] ^ d[511-17] ^ d[511-16] ^ d[511-13] ^ d[511-12] ^ d[511-11] ^ d[511-9] ^ d[511-7] ^ d[511-6] ^ d[511-1] ^ d[511-0] ^ c[31-4] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-16] ^ c[31-20] ^ c[31-23] ^ c[31-26] ^ c[31-29] ^ c[31-30];
                stage_crc512_crc[29] <= d[511-508] ^ d[511-506] ^ d[511-504] ^ d[511-502] ^ d[511-500] ^ d[511-497] ^ d[511-495] ^ d[511-494] ^ d[511-493] ^ d[511-492] ^ d[511-491] ^ d[511-490] ^ d[511-487] ^ d[511-486] ^ d[511-485] ^ d[511-483] ^ d[511-482] ^ d[511-481] ^ d[511-476] ^ d[511-474] ^ d[511-473] ^ d[511-471] ^ d[511-469] ^ d[511-468] ^ d[511-467] ^ d[511-461] ^ d[511-460] ^ d[511-459] ^ d[511-458] ^ d[511-454] ^ d[511-453] ^ d[511-450] ^ d[511-448] ^ d[511-446] ^ d[511-445] ^ d[511-444] ^ d[511-439] ^ d[511-433] ^ d[511-426] ^ d[511-425] ^ d[511-423] ^ d[511-422] ^ d[511-421] ^ d[511-417] ^ d[511-415] ^ d[511-413] ^ d[511-412] ^ d[511-411] ^ d[511-409] ^ d[511-404] ^ d[511-402] ^ d[511-400] ^ d[511-397] ^ d[511-396] ^ d[511-395] ^ d[511-393] ^ d[511-392] ^ d[511-388] ^ d[511-386] ^ d[511-383] ^ d[511-382] ^ d[511-381] ^ d[511-380] ^ d[511-379] ^ d[511-377] ^ d[511-375] ^ d[511-373] ^ d[511-372] ^ d[511-371] ^ d[511-367] ^ d[511-366] ^ d[511-365] ^ d[511-362] ^ d[511-361] ^ d[511-359] ^ d[511-357] ^ d[511-355] ^ d[511-354] ^ d[511-353] ^ d[511-351] ^ d[511-349] ^ d[511-339] ^ d[511-335] ^ d[511-333] ^ d[511-330] ^ d[511-327] ^ d[511-324] ^ d[511-322] ^ d[511-321] ^ d[511-320] ^ d[511-319] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-313] ^ d[511-309] ^ d[511-307] ^ d[511-306] ^ d[511-300] ^ d[511-299] ^ d[511-298] ^ d[511-297] ^ d[511-296] ^ d[511-293] ^ d[511-291] ^ d[511-288] ^ d[511-286] ^ d[511-285] ^ d[511-284] ^ d[511-283] ^ d[511-281] ^ d[511-280] ^ d[511-273] ^ d[511-271] ^ d[511-268] ^ d[511-267] ^ d[511-264] ^ d[511-263] ^ d[511-262] ^ d[511-260] ^ d[511-258] ^ d[511-256] ^ d[511-255] ^ d[511-254] ^ d[511-253] ^ d[511-252] ^ d[511-250] ^ d[511-249] ^ d[511-248] ^ d[511-245] ^ d[511-244] ^ d[511-243] ^ d[511-239] ^ d[511-238] ^ d[511-237] ^ d[511-236] ^ d[511-235] ^ d[511-234] ^ d[511-232] ^ d[511-231] ^ d[511-228] ^ d[511-225] ^ d[511-224] ^ d[511-218] ^ d[511-217] ^ d[511-215] ^ d[511-213] ^ d[511-210] ^ d[511-209] ^ d[511-207] ^ d[511-205] ^ d[511-203] ^ d[511-199] ^ d[511-197] ^ d[511-196] ^ d[511-194] ^ d[511-193] ^ d[511-192] ^ d[511-189] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-182] ^ d[511-174] ^ d[511-172] ^ d[511-171] ^ d[511-166] ^ d[511-164] ^ d[511-161] ^ d[511-160] ^ d[511-159] ^ d[511-155] ^ d[511-153] ^ d[511-152] ^ d[511-150] ^ d[511-149] ^ d[511-146] ^ d[511-143] ^ d[511-139] ^ d[511-137] ^ d[511-136] ^ d[511-133] ^ d[511-132] ^ d[511-130] ^ d[511-128] ^ d[511-127] ^ d[511-124] ^ d[511-123] ^ d[511-121] ^ d[511-119] ^ d[511-118] ^ d[511-110] ^ d[511-108] ^ d[511-107] ^ d[511-102] ^ d[511-99] ^ d[511-98] ^ d[511-97] ^ d[511-96] ^ d[511-94] ^ d[511-89] ^ d[511-88] ^ d[511-85] ^ d[511-84] ^ d[511-83] ^ d[511-80] ^ d[511-79] ^ d[511-75] ^ d[511-72] ^ d[511-70] ^ d[511-68] ^ d[511-67] ^ d[511-64] ^ d[511-59] ^ d[511-58] ^ d[511-57] ^ d[511-55] ^ d[511-53] ^ d[511-52] ^ d[511-51] ^ d[511-44] ^ d[511-39] ^ d[511-38] ^ d[511-37] ^ d[511-36] ^ d[511-35] ^ d[511-32] ^ d[511-31] ^ d[511-30] ^ d[511-26] ^ d[511-24] ^ d[511-18] ^ d[511-17] ^ d[511-16] ^ d[511-14] ^ d[511-13] ^ d[511-9] ^ d[511-8] ^ d[511-7] ^ d[511-6] ^ d[511-2] ^ d[511-1] ^ d[511-0] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-17] ^ c[31-20] ^ c[31-22] ^ c[31-24] ^ c[31-26] ^ c[31-28];
                stage_crc512_crc[28] <= d[511-509] ^ d[511-507] ^ d[511-505] ^ d[511-503] ^ d[511-501] ^ d[511-498] ^ d[511-496] ^ d[511-495] ^ d[511-494] ^ d[511-493] ^ d[511-492] ^ d[511-491] ^ d[511-488] ^ d[511-487] ^ d[511-486] ^ d[511-484] ^ d[511-483] ^ d[511-482] ^ d[511-477] ^ d[511-475] ^ d[511-474] ^ d[511-472] ^ d[511-470] ^ d[511-469] ^ d[511-468] ^ d[511-462] ^ d[511-461] ^ d[511-460] ^ d[511-459] ^ d[511-455] ^ d[511-454] ^ d[511-451] ^ d[511-449] ^ d[511-447] ^ d[511-446] ^ d[511-445] ^ d[511-440] ^ d[511-434] ^ d[511-427] ^ d[511-426] ^ d[511-424] ^ d[511-423] ^ d[511-422] ^ d[511-418] ^ d[511-416] ^ d[511-414] ^ d[511-413] ^ d[511-412] ^ d[511-410] ^ d[511-405] ^ d[511-403] ^ d[511-401] ^ d[511-398] ^ d[511-397] ^ d[511-396] ^ d[511-394] ^ d[511-393] ^ d[511-389] ^ d[511-387] ^ d[511-384] ^ d[511-383] ^ d[511-382] ^ d[511-381] ^ d[511-380] ^ d[511-378] ^ d[511-376] ^ d[511-374] ^ d[511-373] ^ d[511-372] ^ d[511-368] ^ d[511-367] ^ d[511-366] ^ d[511-363] ^ d[511-362] ^ d[511-360] ^ d[511-358] ^ d[511-356] ^ d[511-355] ^ d[511-354] ^ d[511-352] ^ d[511-350] ^ d[511-340] ^ d[511-336] ^ d[511-334] ^ d[511-331] ^ d[511-328] ^ d[511-325] ^ d[511-323] ^ d[511-322] ^ d[511-321] ^ d[511-320] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-310] ^ d[511-308] ^ d[511-307] ^ d[511-301] ^ d[511-300] ^ d[511-299] ^ d[511-298] ^ d[511-297] ^ d[511-294] ^ d[511-292] ^ d[511-289] ^ d[511-287] ^ d[511-286] ^ d[511-285] ^ d[511-284] ^ d[511-282] ^ d[511-281] ^ d[511-274] ^ d[511-272] ^ d[511-269] ^ d[511-268] ^ d[511-265] ^ d[511-264] ^ d[511-263] ^ d[511-261] ^ d[511-259] ^ d[511-257] ^ d[511-256] ^ d[511-255] ^ d[511-254] ^ d[511-253] ^ d[511-251] ^ d[511-250] ^ d[511-249] ^ d[511-246] ^ d[511-245] ^ d[511-244] ^ d[511-240] ^ d[511-239] ^ d[511-238] ^ d[511-237] ^ d[511-236] ^ d[511-235] ^ d[511-233] ^ d[511-232] ^ d[511-229] ^ d[511-226] ^ d[511-225] ^ d[511-219] ^ d[511-218] ^ d[511-216] ^ d[511-214] ^ d[511-211] ^ d[511-210] ^ d[511-208] ^ d[511-206] ^ d[511-204] ^ d[511-200] ^ d[511-198] ^ d[511-197] ^ d[511-195] ^ d[511-194] ^ d[511-193] ^ d[511-190] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-183] ^ d[511-175] ^ d[511-173] ^ d[511-172] ^ d[511-167] ^ d[511-165] ^ d[511-162] ^ d[511-161] ^ d[511-160] ^ d[511-156] ^ d[511-154] ^ d[511-153] ^ d[511-151] ^ d[511-150] ^ d[511-147] ^ d[511-144] ^ d[511-140] ^ d[511-138] ^ d[511-137] ^ d[511-134] ^ d[511-133] ^ d[511-131] ^ d[511-129] ^ d[511-128] ^ d[511-125] ^ d[511-124] ^ d[511-122] ^ d[511-120] ^ d[511-119] ^ d[511-111] ^ d[511-109] ^ d[511-108] ^ d[511-103] ^ d[511-100] ^ d[511-99] ^ d[511-98] ^ d[511-97] ^ d[511-95] ^ d[511-90] ^ d[511-89] ^ d[511-86] ^ d[511-85] ^ d[511-84] ^ d[511-81] ^ d[511-80] ^ d[511-76] ^ d[511-73] ^ d[511-71] ^ d[511-69] ^ d[511-68] ^ d[511-65] ^ d[511-60] ^ d[511-59] ^ d[511-58] ^ d[511-56] ^ d[511-54] ^ d[511-53] ^ d[511-52] ^ d[511-45] ^ d[511-40] ^ d[511-39] ^ d[511-38] ^ d[511-37] ^ d[511-36] ^ d[511-33] ^ d[511-32] ^ d[511-31] ^ d[511-27] ^ d[511-25] ^ d[511-19] ^ d[511-18] ^ d[511-17] ^ d[511-15] ^ d[511-14] ^ d[511-10] ^ d[511-9] ^ d[511-8] ^ d[511-7] ^ d[511-3] ^ d[511-2] ^ d[511-1] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-18] ^ c[31-21] ^ c[31-23] ^ c[31-25] ^ c[31-27] ^ c[31-29];
                stage_crc512_crc[27] <= d[511-511] ^ d[511-507] ^ d[511-504] ^ d[511-501] ^ d[511-500] ^ d[511-499] ^ d[511-497] ^ d[511-496] ^ d[511-491] ^ d[511-490] ^ d[511-487] ^ d[511-486] ^ d[511-485] ^ d[511-484] ^ d[511-482] ^ d[511-481] ^ d[511-480] ^ d[511-479] ^ d[511-478] ^ d[511-477] ^ d[511-475] ^ d[511-473] ^ d[511-472] ^ d[511-471] ^ d[511-469] ^ d[511-468] ^ d[511-465] ^ d[511-464] ^ d[511-463] ^ d[511-460] ^ d[511-458] ^ d[511-456] ^ d[511-455] ^ d[511-449] ^ d[511-447] ^ d[511-446] ^ d[511-444] ^ d[511-441] ^ d[511-437] ^ d[511-436] ^ d[511-435] ^ d[511-434] ^ d[511-433] ^ d[511-428] ^ d[511-427] ^ d[511-425] ^ d[511-423] ^ d[511-422] ^ d[511-418] ^ d[511-417] ^ d[511-416] ^ d[511-415] ^ d[511-413] ^ d[511-412] ^ d[511-411] ^ d[511-409] ^ d[511-408] ^ d[511-407] ^ d[511-406] ^ d[511-405] ^ d[511-402] ^ d[511-400] ^ d[511-397] ^ d[511-396] ^ d[511-395] ^ d[511-394] ^ d[511-393] ^ d[511-392] ^ d[511-391] ^ d[511-387] ^ d[511-386] ^ d[511-385] ^ d[511-384] ^ d[511-383] ^ d[511-382] ^ d[511-379] ^ d[511-378] ^ d[511-377] ^ d[511-376] ^ d[511-375] ^ d[511-373] ^ d[511-372] ^ d[511-367] ^ d[511-366] ^ d[511-364] ^ d[511-362] ^ d[511-361] ^ d[511-358] ^ d[511-356] ^ d[511-355] ^ d[511-351] ^ d[511-349] ^ d[511-348] ^ d[511-347] ^ d[511-345] ^ d[511-344] ^ d[511-342] ^ d[511-339] ^ d[511-338] ^ d[511-334] ^ d[511-333] ^ d[511-332] ^ d[511-329] ^ d[511-328] ^ d[511-327] ^ d[511-326] ^ d[511-324] ^ d[511-323] ^ d[511-320] ^ d[511-319] ^ d[511-316] ^ d[511-312] ^ d[511-311] ^ d[511-310] ^ d[511-308] ^ d[511-305] ^ d[511-303] ^ d[511-301] ^ d[511-297] ^ d[511-296] ^ d[511-294] ^ d[511-293] ^ d[511-292] ^ d[511-285] ^ d[511-282] ^ d[511-279] ^ d[511-277] ^ d[511-276] ^ d[511-275] ^ d[511-274] ^ d[511-270] ^ d[511-268] ^ d[511-266] ^ d[511-262] ^ d[511-261] ^ d[511-260] ^ d[511-259] ^ d[511-258] ^ d[511-256] ^ d[511-254] ^ d[511-251] ^ d[511-250] ^ d[511-248] ^ d[511-247] ^ d[511-246] ^ d[511-245] ^ d[511-243] ^ d[511-241] ^ d[511-240] ^ d[511-239] ^ d[511-238] ^ d[511-236] ^ d[511-233] ^ d[511-228] ^ d[511-224] ^ d[511-220] ^ d[511-219] ^ d[511-217] ^ d[511-216] ^ d[511-215] ^ d[511-214] ^ d[511-211] ^ d[511-210] ^ d[511-208] ^ d[511-205] ^ d[511-203] ^ d[511-202] ^ d[511-197] ^ d[511-196] ^ d[511-195] ^ d[511-193] ^ d[511-192] ^ d[511-190] ^ d[511-189] ^ d[511-187] ^ d[511-186] ^ d[511-184] ^ d[511-183] ^ d[511-182] ^ d[511-176] ^ d[511-174] ^ d[511-173] ^ d[511-172] ^ d[511-171] ^ d[511-170] ^ d[511-169] ^ d[511-168] ^ d[511-167] ^ d[511-163] ^ d[511-158] ^ d[511-157] ^ d[511-156] ^ d[511-154] ^ d[511-152] ^ d[511-149] ^ d[511-148] ^ d[511-145] ^ d[511-144] ^ d[511-143] ^ d[511-141] ^ d[511-139] ^ d[511-138] ^ d[511-137] ^ d[511-136] ^ d[511-130] ^ d[511-129] ^ d[511-128] ^ d[511-127] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-118] ^ d[511-117] ^ d[511-116] ^ d[511-114] ^ d[511-113] ^ d[511-112] ^ d[511-111] ^ d[511-109] ^ d[511-106] ^ d[511-103] ^ d[511-100] ^ d[511-97] ^ d[511-95] ^ d[511-94] ^ d[511-91] ^ d[511-90] ^ d[511-86] ^ d[511-84] ^ d[511-83] ^ d[511-79] ^ d[511-77] ^ d[511-74] ^ d[511-73] ^ d[511-70] ^ d[511-69] ^ d[511-68] ^ d[511-67] ^ d[511-65] ^ d[511-63] ^ d[511-59] ^ d[511-58] ^ d[511-57] ^ d[511-50] ^ d[511-48] ^ d[511-47] ^ d[511-46] ^ d[511-45] ^ d[511-44] ^ d[511-41] ^ d[511-40] ^ d[511-39] ^ d[511-38] ^ d[511-33] ^ d[511-31] ^ d[511-30] ^ d[511-29] ^ d[511-25] ^ d[511-24] ^ d[511-20] ^ d[511-19] ^ d[511-18] ^ d[511-15] ^ d[511-12] ^ d[511-11] ^ d[511-8] ^ d[511-6] ^ d[511-4] ^ d[511-3] ^ d[511-2] ^ d[511-0] ^ c[31-0] ^ c[31-1] ^ c[31-2] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-10] ^ c[31-11] ^ c[31-16] ^ c[31-17] ^ c[31-19] ^ c[31-20] ^ c[31-21] ^ c[31-24] ^ c[31-27] ^ c[31-31];
                stage_crc512_crc[26] <= d[511-511] ^ d[511-510] ^ d[511-507] ^ d[511-506] ^ d[511-505] ^ d[511-498] ^ d[511-497] ^ d[511-495] ^ d[511-494] ^ d[511-493] ^ d[511-490] ^ d[511-489] ^ d[511-487] ^ d[511-485] ^ d[511-478] ^ d[511-477] ^ d[511-474] ^ d[511-473] ^ d[511-469] ^ d[511-468] ^ d[511-466] ^ d[511-462] ^ d[511-459] ^ d[511-458] ^ d[511-457] ^ d[511-456] ^ d[511-452] ^ d[511-449] ^ d[511-447] ^ d[511-445] ^ d[511-444] ^ d[511-442] ^ d[511-438] ^ d[511-435] ^ d[511-433] ^ d[511-429] ^ d[511-428] ^ d[511-426] ^ d[511-423] ^ d[511-422] ^ d[511-417] ^ d[511-413] ^ d[511-410] ^ d[511-406] ^ d[511-405] ^ d[511-404] ^ d[511-403] ^ d[511-401] ^ d[511-400] ^ d[511-399] ^ d[511-397] ^ d[511-395] ^ d[511-394] ^ d[511-391] ^ d[511-390] ^ d[511-385] ^ d[511-384] ^ d[511-383] ^ d[511-381] ^ d[511-380] ^ d[511-379] ^ d[511-377] ^ d[511-373] ^ d[511-372] ^ d[511-369] ^ d[511-367] ^ d[511-366] ^ d[511-365] ^ d[511-358] ^ d[511-356] ^ d[511-353] ^ d[511-352] ^ d[511-350] ^ d[511-347] ^ d[511-346] ^ d[511-344] ^ d[511-343] ^ d[511-342] ^ d[511-341] ^ d[511-340] ^ d[511-338] ^ d[511-337] ^ d[511-330] ^ d[511-329] ^ d[511-325] ^ d[511-324] ^ d[511-322] ^ d[511-319] ^ d[511-318] ^ d[511-315] ^ d[511-313] ^ d[511-311] ^ d[511-310] ^ d[511-306] ^ d[511-305] ^ d[511-304] ^ d[511-303] ^ d[511-300] ^ d[511-299] ^ d[511-296] ^ d[511-293] ^ d[511-292] ^ d[511-290] ^ d[511-288] ^ d[511-287] ^ d[511-280] ^ d[511-279] ^ d[511-278] ^ d[511-275] ^ d[511-274] ^ d[511-273] ^ d[511-271] ^ d[511-268] ^ d[511-267] ^ d[511-265] ^ d[511-264] ^ d[511-263] ^ d[511-262] ^ d[511-260] ^ d[511-251] ^ d[511-249] ^ d[511-247] ^ d[511-246] ^ d[511-244] ^ d[511-243] ^ d[511-242] ^ d[511-241] ^ d[511-240] ^ d[511-239] ^ d[511-230] ^ d[511-229] ^ d[511-228] ^ d[511-227] ^ d[511-226] ^ d[511-225] ^ d[511-224] ^ d[511-221] ^ d[511-220] ^ d[511-218] ^ d[511-217] ^ d[511-215] ^ d[511-214] ^ d[511-211] ^ d[511-210] ^ d[511-208] ^ d[511-207] ^ d[511-206] ^ d[511-204] ^ d[511-202] ^ d[511-201] ^ d[511-199] ^ d[511-196] ^ d[511-192] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-184] ^ d[511-182] ^ d[511-177] ^ d[511-175] ^ d[511-174] ^ d[511-173] ^ d[511-168] ^ d[511-167] ^ d[511-166] ^ d[511-164] ^ d[511-162] ^ d[511-161] ^ d[511-159] ^ d[511-157] ^ d[511-156] ^ d[511-153] ^ d[511-151] ^ d[511-150] ^ d[511-146] ^ d[511-145] ^ d[511-143] ^ d[511-142] ^ d[511-140] ^ d[511-139] ^ d[511-138] ^ d[511-136] ^ d[511-135] ^ d[511-134] ^ d[511-132] ^ d[511-131] ^ d[511-130] ^ d[511-129] ^ d[511-127] ^ d[511-126] ^ d[511-125] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-116] ^ d[511-115] ^ d[511-112] ^ d[511-111] ^ d[511-107] ^ d[511-106] ^ d[511-103] ^ d[511-99] ^ d[511-97] ^ d[511-94] ^ d[511-92] ^ d[511-91] ^ d[511-83] ^ d[511-82] ^ d[511-81] ^ d[511-80] ^ d[511-79] ^ d[511-78] ^ d[511-75] ^ d[511-74] ^ d[511-73] ^ d[511-72] ^ d[511-71] ^ d[511-70] ^ d[511-69] ^ d[511-67] ^ d[511-65] ^ d[511-64] ^ d[511-63] ^ d[511-61] ^ d[511-59] ^ d[511-55] ^ d[511-54] ^ d[511-53] ^ d[511-51] ^ d[511-50] ^ d[511-49] ^ d[511-46] ^ d[511-44] ^ d[511-42] ^ d[511-41] ^ d[511-40] ^ d[511-39] ^ d[511-37] ^ d[511-29] ^ d[511-28] ^ d[511-24] ^ d[511-21] ^ d[511-20] ^ d[511-19] ^ d[511-13] ^ d[511-10] ^ d[511-7] ^ d[511-6] ^ d[511-5] ^ d[511-4] ^ d[511-3] ^ d[511-1] ^ d[511-0] ^ c[31-5] ^ c[31-7] ^ c[31-9] ^ c[31-10] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-17] ^ c[31-18] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-30] ^ c[31-31];
                stage_crc512_crc[25] <= d[511-511] ^ d[511-508] ^ d[511-507] ^ d[511-506] ^ d[511-499] ^ d[511-498] ^ d[511-496] ^ d[511-495] ^ d[511-494] ^ d[511-491] ^ d[511-490] ^ d[511-488] ^ d[511-486] ^ d[511-479] ^ d[511-478] ^ d[511-475] ^ d[511-474] ^ d[511-470] ^ d[511-469] ^ d[511-467] ^ d[511-463] ^ d[511-460] ^ d[511-459] ^ d[511-458] ^ d[511-457] ^ d[511-453] ^ d[511-450] ^ d[511-448] ^ d[511-446] ^ d[511-445] ^ d[511-443] ^ d[511-439] ^ d[511-436] ^ d[511-434] ^ d[511-430] ^ d[511-429] ^ d[511-427] ^ d[511-424] ^ d[511-423] ^ d[511-418] ^ d[511-414] ^ d[511-411] ^ d[511-407] ^ d[511-406] ^ d[511-405] ^ d[511-404] ^ d[511-402] ^ d[511-401] ^ d[511-400] ^ d[511-398] ^ d[511-396] ^ d[511-395] ^ d[511-392] ^ d[511-391] ^ d[511-386] ^ d[511-385] ^ d[511-384] ^ d[511-382] ^ d[511-381] ^ d[511-380] ^ d[511-378] ^ d[511-374] ^ d[511-373] ^ d[511-370] ^ d[511-368] ^ d[511-367] ^ d[511-366] ^ d[511-359] ^ d[511-357] ^ d[511-354] ^ d[511-353] ^ d[511-351] ^ d[511-348] ^ d[511-347] ^ d[511-345] ^ d[511-344] ^ d[511-343] ^ d[511-342] ^ d[511-341] ^ d[511-339] ^ d[511-338] ^ d[511-331] ^ d[511-330] ^ d[511-326] ^ d[511-325] ^ d[511-323] ^ d[511-320] ^ d[511-319] ^ d[511-316] ^ d[511-314] ^ d[511-312] ^ d[511-311] ^ d[511-307] ^ d[511-306] ^ d[511-305] ^ d[511-304] ^ d[511-301] ^ d[511-300] ^ d[511-297] ^ d[511-294] ^ d[511-293] ^ d[511-291] ^ d[511-289] ^ d[511-288] ^ d[511-281] ^ d[511-280] ^ d[511-279] ^ d[511-276] ^ d[511-275] ^ d[511-274] ^ d[511-272] ^ d[511-269] ^ d[511-268] ^ d[511-266] ^ d[511-265] ^ d[511-264] ^ d[511-263] ^ d[511-261] ^ d[511-252] ^ d[511-250] ^ d[511-248] ^ d[511-247] ^ d[511-245] ^ d[511-244] ^ d[511-243] ^ d[511-242] ^ d[511-241] ^ d[511-240] ^ d[511-231] ^ d[511-230] ^ d[511-229] ^ d[511-228] ^ d[511-227] ^ d[511-226] ^ d[511-225] ^ d[511-222] ^ d[511-221] ^ d[511-219] ^ d[511-218] ^ d[511-216] ^ d[511-215] ^ d[511-212] ^ d[511-211] ^ d[511-209] ^ d[511-208] ^ d[511-207] ^ d[511-205] ^ d[511-203] ^ d[511-202] ^ d[511-200] ^ d[511-197] ^ d[511-193] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-183] ^ d[511-178] ^ d[511-176] ^ d[511-175] ^ d[511-174] ^ d[511-169] ^ d[511-168] ^ d[511-167] ^ d[511-165] ^ d[511-163] ^ d[511-162] ^ d[511-160] ^ d[511-158] ^ d[511-157] ^ d[511-154] ^ d[511-152] ^ d[511-151] ^ d[511-147] ^ d[511-146] ^ d[511-144] ^ d[511-143] ^ d[511-141] ^ d[511-140] ^ d[511-139] ^ d[511-137] ^ d[511-136] ^ d[511-135] ^ d[511-133] ^ d[511-132] ^ d[511-131] ^ d[511-130] ^ d[511-128] ^ d[511-127] ^ d[511-126] ^ d[511-124] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-117] ^ d[511-116] ^ d[511-113] ^ d[511-112] ^ d[511-108] ^ d[511-107] ^ d[511-104] ^ d[511-100] ^ d[511-98] ^ d[511-95] ^ d[511-93] ^ d[511-92] ^ d[511-84] ^ d[511-83] ^ d[511-82] ^ d[511-81] ^ d[511-80] ^ d[511-79] ^ d[511-76] ^ d[511-75] ^ d[511-74] ^ d[511-73] ^ d[511-72] ^ d[511-71] ^ d[511-70] ^ d[511-68] ^ d[511-66] ^ d[511-65] ^ d[511-64] ^ d[511-62] ^ d[511-60] ^ d[511-56] ^ d[511-55] ^ d[511-54] ^ d[511-52] ^ d[511-51] ^ d[511-50] ^ d[511-47] ^ d[511-45] ^ d[511-43] ^ d[511-42] ^ d[511-41] ^ d[511-40] ^ d[511-38] ^ d[511-30] ^ d[511-29] ^ d[511-25] ^ d[511-22] ^ d[511-21] ^ d[511-20] ^ d[511-14] ^ d[511-11] ^ d[511-8] ^ d[511-7] ^ d[511-6] ^ d[511-5] ^ d[511-4] ^ d[511-2] ^ d[511-1] ^ c[31-6] ^ c[31-8] ^ c[31-10] ^ c[31-11] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-18] ^ c[31-19] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-31];
                stage_crc512_crc[24] <= d[511-511] ^ d[511-510] ^ d[511-509] ^ d[511-506] ^ d[511-502] ^ d[511-501] ^ d[511-499] ^ d[511-497] ^ d[511-496] ^ d[511-494] ^ d[511-493] ^ d[511-490] ^ d[511-488] ^ d[511-487] ^ d[511-486] ^ d[511-483] ^ d[511-482] ^ d[511-481] ^ d[511-477] ^ d[511-475] ^ d[511-472] ^ d[511-471] ^ d[511-465] ^ d[511-462] ^ d[511-460] ^ d[511-459] ^ d[511-454] ^ d[511-452] ^ d[511-451] ^ d[511-450] ^ d[511-448] ^ d[511-447] ^ d[511-446] ^ d[511-440] ^ d[511-436] ^ d[511-435] ^ d[511-434] ^ d[511-433] ^ d[511-431] ^ d[511-430] ^ d[511-428] ^ d[511-425] ^ d[511-422] ^ d[511-418] ^ d[511-416] ^ d[511-415] ^ d[511-414] ^ d[511-409] ^ d[511-406] ^ d[511-404] ^ d[511-403] ^ d[511-402] ^ d[511-401] ^ d[511-400] ^ d[511-398] ^ d[511-397] ^ d[511-391] ^ d[511-390] ^ d[511-388] ^ d[511-385] ^ d[511-383] ^ d[511-382] ^ d[511-379] ^ d[511-378] ^ d[511-376] ^ d[511-375] ^ d[511-372] ^ d[511-371] ^ d[511-367] ^ d[511-366] ^ d[511-363] ^ d[511-362] ^ d[511-360] ^ d[511-359] ^ d[511-357] ^ d[511-355] ^ d[511-354] ^ d[511-353] ^ d[511-352] ^ d[511-347] ^ d[511-346] ^ d[511-343] ^ d[511-341] ^ d[511-340] ^ d[511-338] ^ d[511-337] ^ d[511-335] ^ d[511-334] ^ d[511-333] ^ d[511-332] ^ d[511-331] ^ d[511-328] ^ d[511-326] ^ d[511-324] ^ d[511-322] ^ d[511-319] ^ d[511-318] ^ d[511-313] ^ d[511-310] ^ d[511-309] ^ d[511-308] ^ d[511-307] ^ d[511-306] ^ d[511-303] ^ d[511-301] ^ d[511-300] ^ d[511-299] ^ d[511-297] ^ d[511-296] ^ d[511-289] ^ d[511-288] ^ d[511-287] ^ d[511-286] ^ d[511-283] ^ d[511-282] ^ d[511-281] ^ d[511-280] ^ d[511-279] ^ d[511-275] ^ d[511-274] ^ d[511-270] ^ d[511-268] ^ d[511-267] ^ d[511-266] ^ d[511-262] ^ d[511-261] ^ d[511-259] ^ d[511-257] ^ d[511-255] ^ d[511-253] ^ d[511-252] ^ d[511-251] ^ d[511-249] ^ d[511-246] ^ d[511-245] ^ d[511-244] ^ d[511-242] ^ d[511-241] ^ d[511-237] ^ d[511-234] ^ d[511-232] ^ d[511-231] ^ d[511-229] ^ d[511-224] ^ d[511-223] ^ d[511-222] ^ d[511-220] ^ d[511-219] ^ d[511-217] ^ d[511-214] ^ d[511-213] ^ d[511-207] ^ d[511-206] ^ d[511-204] ^ d[511-202] ^ d[511-199] ^ d[511-197] ^ d[511-193] ^ d[511-192] ^ d[511-191] ^ d[511-190] ^ d[511-189] ^ d[511-187] ^ d[511-184] ^ d[511-183] ^ d[511-182] ^ d[511-179] ^ d[511-177] ^ d[511-176] ^ d[511-175] ^ d[511-172] ^ d[511-171] ^ d[511-168] ^ d[511-167] ^ d[511-164] ^ d[511-163] ^ d[511-162] ^ d[511-159] ^ d[511-156] ^ d[511-153] ^ d[511-152] ^ d[511-151] ^ d[511-149] ^ d[511-148] ^ d[511-147] ^ d[511-145] ^ d[511-143] ^ d[511-142] ^ d[511-141] ^ d[511-140] ^ d[511-138] ^ d[511-135] ^ d[511-133] ^ d[511-131] ^ d[511-129] ^ d[511-126] ^ d[511-124] ^ d[511-122] ^ d[511-119] ^ d[511-116] ^ d[511-111] ^ d[511-110] ^ d[511-109] ^ d[511-108] ^ d[511-106] ^ d[511-105] ^ d[511-104] ^ d[511-103] ^ d[511-98] ^ d[511-97] ^ d[511-95] ^ d[511-93] ^ d[511-87] ^ d[511-80] ^ d[511-79] ^ d[511-77] ^ d[511-76] ^ d[511-75] ^ d[511-74] ^ d[511-71] ^ d[511-69] ^ d[511-68] ^ d[511-60] ^ d[511-58] ^ d[511-57] ^ d[511-56] ^ d[511-54] ^ d[511-52] ^ d[511-51] ^ d[511-50] ^ d[511-47] ^ d[511-46] ^ d[511-45] ^ d[511-43] ^ d[511-42] ^ d[511-41] ^ d[511-39] ^ d[511-37] ^ d[511-34] ^ d[511-32] ^ d[511-29] ^ d[511-28] ^ d[511-25] ^ d[511-24] ^ d[511-23] ^ d[511-22] ^ d[511-21] ^ d[511-16] ^ d[511-15] ^ d[511-10] ^ d[511-8] ^ d[511-7] ^ d[511-5] ^ d[511-3] ^ d[511-2] ^ d[511-0] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-10] ^ c[31-13] ^ c[31-14] ^ c[31-16] ^ c[31-17] ^ c[31-19] ^ c[31-21] ^ c[31-22] ^ c[31-26] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc512_crc[23] <= d[511-508] ^ d[511-506] ^ d[511-503] ^ d[511-501] ^ d[511-498] ^ d[511-497] ^ d[511-493] ^ d[511-492] ^ d[511-490] ^ d[511-487] ^ d[511-486] ^ d[511-484] ^ d[511-481] ^ d[511-480] ^ d[511-479] ^ d[511-478] ^ d[511-477] ^ d[511-473] ^ d[511-470] ^ d[511-468] ^ d[511-466] ^ d[511-465] ^ d[511-464] ^ d[511-463] ^ d[511-462] ^ d[511-460] ^ d[511-458] ^ d[511-455] ^ d[511-453] ^ d[511-451] ^ d[511-450] ^ d[511-447] ^ d[511-444] ^ d[511-441] ^ d[511-435] ^ d[511-433] ^ d[511-432] ^ d[511-431] ^ d[511-429] ^ d[511-426] ^ d[511-424] ^ d[511-423] ^ d[511-422] ^ d[511-418] ^ d[511-417] ^ d[511-415] ^ d[511-414] ^ d[511-412] ^ d[511-410] ^ d[511-409] ^ d[511-408] ^ d[511-403] ^ d[511-402] ^ d[511-401] ^ d[511-400] ^ d[511-396] ^ d[511-393] ^ d[511-390] ^ d[511-389] ^ d[511-388] ^ d[511-387] ^ d[511-384] ^ d[511-383] ^ d[511-381] ^ d[511-380] ^ d[511-379] ^ d[511-378] ^ d[511-377] ^ d[511-374] ^ d[511-373] ^ d[511-369] ^ d[511-367] ^ d[511-366] ^ d[511-364] ^ d[511-362] ^ d[511-361] ^ d[511-360] ^ d[511-359] ^ d[511-357] ^ d[511-356] ^ d[511-355] ^ d[511-354] ^ d[511-349] ^ d[511-345] ^ d[511-337] ^ d[511-336] ^ d[511-332] ^ d[511-329] ^ d[511-328] ^ d[511-325] ^ d[511-323] ^ d[511-322] ^ d[511-321] ^ d[511-318] ^ d[511-317] ^ d[511-315] ^ d[511-314] ^ d[511-312] ^ d[511-311] ^ d[511-308] ^ d[511-307] ^ d[511-305] ^ d[511-304] ^ d[511-303] ^ d[511-301] ^ d[511-299] ^ d[511-296] ^ d[511-295] ^ d[511-294] ^ d[511-292] ^ d[511-289] ^ d[511-286] ^ d[511-284] ^ d[511-282] ^ d[511-281] ^ d[511-280] ^ d[511-279] ^ d[511-277] ^ d[511-275] ^ d[511-274] ^ d[511-273] ^ d[511-271] ^ d[511-267] ^ d[511-265] ^ d[511-264] ^ d[511-263] ^ d[511-262] ^ d[511-261] ^ d[511-260] ^ d[511-259] ^ d[511-258] ^ d[511-257] ^ d[511-256] ^ d[511-255] ^ d[511-254] ^ d[511-253] ^ d[511-250] ^ d[511-248] ^ d[511-247] ^ d[511-246] ^ d[511-245] ^ d[511-242] ^ d[511-238] ^ d[511-237] ^ d[511-235] ^ d[511-234] ^ d[511-233] ^ d[511-232] ^ d[511-228] ^ d[511-227] ^ d[511-226] ^ d[511-225] ^ d[511-223] ^ d[511-221] ^ d[511-220] ^ d[511-218] ^ d[511-216] ^ d[511-215] ^ d[511-212] ^ d[511-210] ^ d[511-209] ^ d[511-205] ^ d[511-202] ^ d[511-201] ^ d[511-200] ^ d[511-199] ^ d[511-197] ^ d[511-186] ^ d[511-185] ^ d[511-184] ^ d[511-182] ^ d[511-180] ^ d[511-178] ^ d[511-177] ^ d[511-176] ^ d[511-173] ^ d[511-171] ^ d[511-170] ^ d[511-168] ^ d[511-167] ^ d[511-166] ^ d[511-165] ^ d[511-164] ^ d[511-163] ^ d[511-162] ^ d[511-161] ^ d[511-160] ^ d[511-158] ^ d[511-157] ^ d[511-156] ^ d[511-155] ^ d[511-154] ^ d[511-153] ^ d[511-152] ^ d[511-151] ^ d[511-150] ^ d[511-148] ^ d[511-146] ^ d[511-142] ^ d[511-141] ^ d[511-139] ^ d[511-137] ^ d[511-135] ^ d[511-130] ^ d[511-128] ^ d[511-126] ^ d[511-120] ^ d[511-119] ^ d[511-118] ^ d[511-116] ^ d[511-114] ^ d[511-113] ^ d[511-112] ^ d[511-109] ^ d[511-107] ^ d[511-105] ^ d[511-103] ^ d[511-101] ^ d[511-97] ^ d[511-95] ^ d[511-88] ^ d[511-87] ^ d[511-85] ^ d[511-84] ^ d[511-83] ^ d[511-82] ^ d[511-80] ^ d[511-79] ^ d[511-78] ^ d[511-77] ^ d[511-76] ^ d[511-75] ^ d[511-73] ^ d[511-70] ^ d[511-69] ^ d[511-68] ^ d[511-67] ^ d[511-66] ^ d[511-65] ^ d[511-63] ^ d[511-60] ^ d[511-59] ^ d[511-57] ^ d[511-54] ^ d[511-52] ^ d[511-51] ^ d[511-50] ^ d[511-46] ^ d[511-45] ^ d[511-43] ^ d[511-42] ^ d[511-40] ^ d[511-38] ^ d[511-37] ^ d[511-35] ^ d[511-34] ^ d[511-33] ^ d[511-32] ^ d[511-31] ^ d[511-28] ^ d[511-23] ^ d[511-22] ^ d[511-17] ^ d[511-12] ^ d[511-11] ^ d[511-10] ^ d[511-8] ^ d[511-4] ^ d[511-3] ^ d[511-1] ^ d[511-0] ^ c[31-0] ^ c[31-1] ^ c[31-4] ^ c[31-6] ^ c[31-7] ^ c[31-10] ^ c[31-12] ^ c[31-13] ^ c[31-17] ^ c[31-18] ^ c[31-21] ^ c[31-23] ^ c[31-26] ^ c[31-28];
                stage_crc512_crc[22] <= d[511-509] ^ d[511-507] ^ d[511-504] ^ d[511-502] ^ d[511-499] ^ d[511-498] ^ d[511-494] ^ d[511-493] ^ d[511-491] ^ d[511-488] ^ d[511-487] ^ d[511-485] ^ d[511-482] ^ d[511-481] ^ d[511-480] ^ d[511-479] ^ d[511-478] ^ d[511-474] ^ d[511-471] ^ d[511-469] ^ d[511-467] ^ d[511-466] ^ d[511-465] ^ d[511-464] ^ d[511-463] ^ d[511-461] ^ d[511-459] ^ d[511-456] ^ d[511-454] ^ d[511-452] ^ d[511-451] ^ d[511-448] ^ d[511-445] ^ d[511-442] ^ d[511-436] ^ d[511-434] ^ d[511-433] ^ d[511-432] ^ d[511-430] ^ d[511-427] ^ d[511-425] ^ d[511-424] ^ d[511-423] ^ d[511-419] ^ d[511-418] ^ d[511-416] ^ d[511-415] ^ d[511-413] ^ d[511-411] ^ d[511-410] ^ d[511-409] ^ d[511-404] ^ d[511-403] ^ d[511-402] ^ d[511-401] ^ d[511-397] ^ d[511-394] ^ d[511-391] ^ d[511-390] ^ d[511-389] ^ d[511-388] ^ d[511-385] ^ d[511-384] ^ d[511-382] ^ d[511-381] ^ d[511-380] ^ d[511-379] ^ d[511-378] ^ d[511-375] ^ d[511-374] ^ d[511-370] ^ d[511-368] ^ d[511-367] ^ d[511-365] ^ d[511-363] ^ d[511-362] ^ d[511-361] ^ d[511-360] ^ d[511-358] ^ d[511-357] ^ d[511-356] ^ d[511-355] ^ d[511-350] ^ d[511-346] ^ d[511-338] ^ d[511-337] ^ d[511-333] ^ d[511-330] ^ d[511-329] ^ d[511-326] ^ d[511-324] ^ d[511-323] ^ d[511-322] ^ d[511-319] ^ d[511-318] ^ d[511-316] ^ d[511-315] ^ d[511-313] ^ d[511-312] ^ d[511-309] ^ d[511-308] ^ d[511-306] ^ d[511-305] ^ d[511-304] ^ d[511-302] ^ d[511-300] ^ d[511-297] ^ d[511-296] ^ d[511-295] ^ d[511-293] ^ d[511-290] ^ d[511-287] ^ d[511-285] ^ d[511-283] ^ d[511-282] ^ d[511-281] ^ d[511-280] ^ d[511-278] ^ d[511-276] ^ d[511-275] ^ d[511-274] ^ d[511-272] ^ d[511-268] ^ d[511-266] ^ d[511-265] ^ d[511-264] ^ d[511-263] ^ d[511-262] ^ d[511-261] ^ d[511-260] ^ d[511-259] ^ d[511-258] ^ d[511-257] ^ d[511-256] ^ d[511-255] ^ d[511-254] ^ d[511-251] ^ d[511-249] ^ d[511-248] ^ d[511-247] ^ d[511-246] ^ d[511-243] ^ d[511-239] ^ d[511-238] ^ d[511-236] ^ d[511-235] ^ d[511-234] ^ d[511-233] ^ d[511-229] ^ d[511-228] ^ d[511-227] ^ d[511-226] ^ d[511-224] ^ d[511-222] ^ d[511-221] ^ d[511-219] ^ d[511-217] ^ d[511-216] ^ d[511-213] ^ d[511-211] ^ d[511-210] ^ d[511-206] ^ d[511-203] ^ d[511-202] ^ d[511-201] ^ d[511-200] ^ d[511-198] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-183] ^ d[511-181] ^ d[511-179] ^ d[511-178] ^ d[511-177] ^ d[511-174] ^ d[511-172] ^ d[511-171] ^ d[511-169] ^ d[511-168] ^ d[511-167] ^ d[511-166] ^ d[511-165] ^ d[511-164] ^ d[511-163] ^ d[511-162] ^ d[511-161] ^ d[511-159] ^ d[511-158] ^ d[511-157] ^ d[511-156] ^ d[511-155] ^ d[511-154] ^ d[511-153] ^ d[511-152] ^ d[511-151] ^ d[511-149] ^ d[511-147] ^ d[511-143] ^ d[511-142] ^ d[511-140] ^ d[511-138] ^ d[511-136] ^ d[511-131] ^ d[511-129] ^ d[511-127] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-117] ^ d[511-115] ^ d[511-114] ^ d[511-113] ^ d[511-110] ^ d[511-108] ^ d[511-106] ^ d[511-104] ^ d[511-102] ^ d[511-98] ^ d[511-96] ^ d[511-89] ^ d[511-88] ^ d[511-86] ^ d[511-85] ^ d[511-84] ^ d[511-83] ^ d[511-81] ^ d[511-80] ^ d[511-79] ^ d[511-78] ^ d[511-77] ^ d[511-76] ^ d[511-74] ^ d[511-71] ^ d[511-70] ^ d[511-69] ^ d[511-68] ^ d[511-67] ^ d[511-66] ^ d[511-64] ^ d[511-61] ^ d[511-60] ^ d[511-58] ^ d[511-55] ^ d[511-53] ^ d[511-52] ^ d[511-51] ^ d[511-47] ^ d[511-46] ^ d[511-44] ^ d[511-43] ^ d[511-41] ^ d[511-39] ^ d[511-38] ^ d[511-36] ^ d[511-35] ^ d[511-34] ^ d[511-33] ^ d[511-32] ^ d[511-29] ^ d[511-24] ^ d[511-23] ^ d[511-18] ^ d[511-13] ^ d[511-12] ^ d[511-11] ^ d[511-9] ^ d[511-5] ^ d[511-4] ^ d[511-2] ^ d[511-1] ^ c[31-0] ^ c[31-1] ^ c[31-2] ^ c[31-5] ^ c[31-7] ^ c[31-8] ^ c[31-11] ^ c[31-13] ^ c[31-14] ^ c[31-18] ^ c[31-19] ^ c[31-22] ^ c[31-24] ^ c[31-27] ^ c[31-29];
                stage_crc512_crc[21] <= d[511-511] ^ d[511-507] ^ d[511-506] ^ d[511-505] ^ d[511-503] ^ d[511-502] ^ d[511-501] ^ d[511-499] ^ d[511-493] ^ d[511-491] ^ d[511-490] ^ d[511-477] ^ d[511-476] ^ d[511-475] ^ d[511-467] ^ d[511-466] ^ d[511-461] ^ d[511-460] ^ d[511-458] ^ d[511-457] ^ d[511-455] ^ d[511-453] ^ d[511-450] ^ d[511-448] ^ d[511-446] ^ d[511-444] ^ d[511-443] ^ d[511-436] ^ d[511-435] ^ d[511-431] ^ d[511-428] ^ d[511-426] ^ d[511-425] ^ d[511-422] ^ d[511-420] ^ d[511-418] ^ d[511-417] ^ d[511-411] ^ d[511-410] ^ d[511-409] ^ d[511-408] ^ d[511-407] ^ d[511-403] ^ d[511-402] ^ d[511-400] ^ d[511-399] ^ d[511-396] ^ d[511-395] ^ d[511-393] ^ d[511-389] ^ d[511-388] ^ d[511-387] ^ d[511-385] ^ d[511-383] ^ d[511-382] ^ d[511-380] ^ d[511-379] ^ d[511-378] ^ d[511-375] ^ d[511-374] ^ d[511-372] ^ d[511-371] ^ d[511-364] ^ d[511-361] ^ d[511-356] ^ d[511-353] ^ d[511-351] ^ d[511-349] ^ d[511-348] ^ d[511-345] ^ d[511-344] ^ d[511-342] ^ d[511-341] ^ d[511-337] ^ d[511-335] ^ d[511-333] ^ d[511-331] ^ d[511-330] ^ d[511-328] ^ d[511-325] ^ d[511-324] ^ d[511-323] ^ d[511-322] ^ d[511-321] ^ d[511-318] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-313] ^ d[511-312] ^ d[511-307] ^ d[511-306] ^ d[511-302] ^ d[511-301] ^ d[511-300] ^ d[511-299] ^ d[511-295] ^ d[511-292] ^ d[511-291] ^ d[511-290] ^ d[511-287] ^ d[511-284] ^ d[511-282] ^ d[511-281] ^ d[511-275] ^ d[511-274] ^ d[511-268] ^ d[511-267] ^ d[511-266] ^ d[511-263] ^ d[511-262] ^ d[511-260] ^ d[511-258] ^ d[511-256] ^ d[511-250] ^ d[511-249] ^ d[511-247] ^ d[511-244] ^ d[511-243] ^ d[511-240] ^ d[511-239] ^ d[511-236] ^ d[511-235] ^ d[511-229] ^ d[511-226] ^ d[511-225] ^ d[511-224] ^ d[511-223] ^ d[511-222] ^ d[511-220] ^ d[511-218] ^ d[511-217] ^ d[511-216] ^ d[511-211] ^ d[511-210] ^ d[511-209] ^ d[511-208] ^ d[511-204] ^ d[511-198] ^ d[511-197] ^ d[511-194] ^ d[511-193] ^ d[511-192] ^ d[511-191] ^ d[511-190] ^ d[511-187] ^ d[511-184] ^ d[511-183] ^ d[511-180] ^ d[511-179] ^ d[511-178] ^ d[511-175] ^ d[511-173] ^ d[511-171] ^ d[511-168] ^ d[511-165] ^ d[511-164] ^ d[511-163] ^ d[511-161] ^ d[511-160] ^ d[511-159] ^ d[511-157] ^ d[511-154] ^ d[511-153] ^ d[511-152] ^ d[511-151] ^ d[511-150] ^ d[511-149] ^ d[511-148] ^ d[511-141] ^ d[511-139] ^ d[511-136] ^ d[511-135] ^ d[511-134] ^ d[511-130] ^ d[511-127] ^ d[511-126] ^ d[511-125] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-117] ^ d[511-115] ^ d[511-113] ^ d[511-110] ^ d[511-109] ^ d[511-107] ^ d[511-106] ^ d[511-105] ^ d[511-104] ^ d[511-101] ^ d[511-98] ^ d[511-96] ^ d[511-95] ^ d[511-94] ^ d[511-90] ^ d[511-89] ^ d[511-86] ^ d[511-83] ^ d[511-80] ^ d[511-78] ^ d[511-77] ^ d[511-75] ^ d[511-73] ^ d[511-71] ^ d[511-70] ^ d[511-69] ^ d[511-66] ^ d[511-63] ^ d[511-62] ^ d[511-60] ^ d[511-59] ^ d[511-58] ^ d[511-56] ^ d[511-55] ^ d[511-52] ^ d[511-50] ^ d[511-42] ^ d[511-40] ^ d[511-39] ^ d[511-36] ^ d[511-35] ^ d[511-33] ^ d[511-32] ^ d[511-31] ^ d[511-29] ^ d[511-28] ^ d[511-26] ^ d[511-19] ^ d[511-16] ^ d[511-14] ^ d[511-13] ^ d[511-9] ^ d[511-5] ^ d[511-3] ^ d[511-2] ^ d[511-0] ^ c[31-10] ^ c[31-11] ^ c[31-13] ^ c[31-19] ^ c[31-21] ^ c[31-22] ^ c[31-23] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-31];
                stage_crc512_crc[20] <= d[511-511] ^ d[511-510] ^ d[511-504] ^ d[511-503] ^ d[511-501] ^ d[511-495] ^ d[511-493] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-486] ^ d[511-483] ^ d[511-482] ^ d[511-481] ^ d[511-480] ^ d[511-479] ^ d[511-478] ^ d[511-472] ^ d[511-470] ^ d[511-467] ^ d[511-465] ^ d[511-464] ^ d[511-459] ^ d[511-456] ^ d[511-454] ^ d[511-452] ^ d[511-451] ^ d[511-450] ^ d[511-448] ^ d[511-447] ^ d[511-445] ^ d[511-434] ^ d[511-433] ^ d[511-432] ^ d[511-429] ^ d[511-427] ^ d[511-426] ^ d[511-424] ^ d[511-423] ^ d[511-422] ^ d[511-421] ^ d[511-416] ^ d[511-414] ^ d[511-411] ^ d[511-410] ^ d[511-407] ^ d[511-405] ^ d[511-403] ^ d[511-401] ^ d[511-399] ^ d[511-398] ^ d[511-397] ^ d[511-394] ^ d[511-393] ^ d[511-392] ^ d[511-391] ^ d[511-389] ^ d[511-387] ^ d[511-384] ^ d[511-383] ^ d[511-380] ^ d[511-379] ^ d[511-378] ^ d[511-375] ^ d[511-374] ^ d[511-373] ^ d[511-369] ^ d[511-368] ^ d[511-366] ^ d[511-365] ^ d[511-363] ^ d[511-359] ^ d[511-358] ^ d[511-354] ^ d[511-353] ^ d[511-352] ^ d[511-350] ^ d[511-348] ^ d[511-347] ^ d[511-346] ^ d[511-344] ^ d[511-343] ^ d[511-341] ^ d[511-339] ^ d[511-337] ^ d[511-336] ^ d[511-335] ^ d[511-333] ^ d[511-332] ^ d[511-331] ^ d[511-329] ^ d[511-328] ^ d[511-327] ^ d[511-326] ^ d[511-325] ^ d[511-324] ^ d[511-323] ^ d[511-321] ^ d[511-320] ^ d[511-318] ^ d[511-316] ^ d[511-314] ^ d[511-313] ^ d[511-312] ^ d[511-310] ^ d[511-309] ^ d[511-308] ^ d[511-307] ^ d[511-305] ^ d[511-301] ^ d[511-299] ^ d[511-298] ^ d[511-297] ^ d[511-295] ^ d[511-294] ^ d[511-293] ^ d[511-291] ^ d[511-290] ^ d[511-287] ^ d[511-286] ^ d[511-285] ^ d[511-282] ^ d[511-279] ^ d[511-277] ^ d[511-275] ^ d[511-274] ^ d[511-273] ^ d[511-267] ^ d[511-265] ^ d[511-263] ^ d[511-255] ^ d[511-252] ^ d[511-251] ^ d[511-250] ^ d[511-245] ^ d[511-244] ^ d[511-243] ^ d[511-241] ^ d[511-240] ^ d[511-236] ^ d[511-234] ^ d[511-228] ^ d[511-225] ^ d[511-223] ^ d[511-221] ^ d[511-219] ^ d[511-218] ^ d[511-217] ^ d[511-216] ^ d[511-214] ^ d[511-211] ^ d[511-208] ^ d[511-207] ^ d[511-205] ^ d[511-203] ^ d[511-202] ^ d[511-201] ^ d[511-197] ^ d[511-195] ^ d[511-190] ^ d[511-186] ^ d[511-185] ^ d[511-184] ^ d[511-183] ^ d[511-182] ^ d[511-181] ^ d[511-180] ^ d[511-179] ^ d[511-176] ^ d[511-174] ^ d[511-171] ^ d[511-170] ^ d[511-167] ^ d[511-165] ^ d[511-164] ^ d[511-160] ^ d[511-156] ^ d[511-154] ^ d[511-153] ^ d[511-152] ^ d[511-150] ^ d[511-144] ^ d[511-143] ^ d[511-142] ^ d[511-140] ^ d[511-134] ^ d[511-132] ^ d[511-131] ^ d[511-125] ^ d[511-124] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-117] ^ d[511-113] ^ d[511-108] ^ d[511-107] ^ d[511-105] ^ d[511-104] ^ d[511-103] ^ d[511-102] ^ d[511-101] ^ d[511-98] ^ d[511-94] ^ d[511-91] ^ d[511-90] ^ d[511-85] ^ d[511-83] ^ d[511-82] ^ d[511-78] ^ d[511-76] ^ d[511-74] ^ d[511-73] ^ d[511-71] ^ d[511-70] ^ d[511-68] ^ d[511-66] ^ d[511-65] ^ d[511-64] ^ d[511-59] ^ d[511-58] ^ d[511-57] ^ d[511-56] ^ d[511-55] ^ d[511-54] ^ d[511-51] ^ d[511-50] ^ d[511-48] ^ d[511-47] ^ d[511-45] ^ d[511-44] ^ d[511-43] ^ d[511-41] ^ d[511-40] ^ d[511-36] ^ d[511-33] ^ d[511-31] ^ d[511-28] ^ d[511-27] ^ d[511-26] ^ d[511-25] ^ d[511-24] ^ d[511-20] ^ d[511-17] ^ d[511-16] ^ d[511-15] ^ d[511-14] ^ d[511-12] ^ d[511-9] ^ d[511-4] ^ d[511-3] ^ d[511-1] ^ d[511-0] ^ c[31-0] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-6] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-13] ^ c[31-15] ^ c[31-21] ^ c[31-23] ^ c[31-24] ^ c[31-30] ^ c[31-31];
                stage_crc512_crc[19] <= d[511-510] ^ d[511-508] ^ d[511-507] ^ d[511-506] ^ d[511-505] ^ d[511-504] ^ d[511-501] ^ d[511-500] ^ d[511-496] ^ d[511-495] ^ d[511-493] ^ d[511-492] ^ d[511-488] ^ d[511-487] ^ d[511-486] ^ d[511-484] ^ d[511-477] ^ d[511-476] ^ d[511-473] ^ d[511-472] ^ d[511-471] ^ d[511-470] ^ d[511-466] ^ d[511-464] ^ d[511-462] ^ d[511-461] ^ d[511-460] ^ d[511-458] ^ d[511-457] ^ d[511-455] ^ d[511-453] ^ d[511-451] ^ d[511-450] ^ d[511-446] ^ d[511-444] ^ d[511-437] ^ d[511-436] ^ d[511-435] ^ d[511-430] ^ d[511-428] ^ d[511-427] ^ d[511-425] ^ d[511-423] ^ d[511-419] ^ d[511-418] ^ d[511-417] ^ d[511-416] ^ d[511-415] ^ d[511-414] ^ d[511-411] ^ d[511-409] ^ d[511-407] ^ d[511-406] ^ d[511-405] ^ d[511-402] ^ d[511-396] ^ d[511-395] ^ d[511-394] ^ d[511-391] ^ d[511-387] ^ d[511-386] ^ d[511-385] ^ d[511-384] ^ d[511-380] ^ d[511-379] ^ d[511-378] ^ d[511-375] ^ d[511-372] ^ d[511-370] ^ d[511-368] ^ d[511-367] ^ d[511-364] ^ d[511-363] ^ d[511-362] ^ d[511-360] ^ d[511-358] ^ d[511-357] ^ d[511-355] ^ d[511-354] ^ d[511-351] ^ d[511-341] ^ d[511-340] ^ d[511-339] ^ d[511-336] ^ d[511-335] ^ d[511-332] ^ d[511-330] ^ d[511-329] ^ d[511-326] ^ d[511-325] ^ d[511-324] ^ d[511-320] ^ d[511-318] ^ d[511-314] ^ d[511-313] ^ d[511-312] ^ d[511-311] ^ d[511-308] ^ d[511-306] ^ d[511-305] ^ d[511-303] ^ d[511-297] ^ d[511-291] ^ d[511-290] ^ d[511-280] ^ d[511-279] ^ d[511-278] ^ d[511-277] ^ d[511-275] ^ d[511-273] ^ d[511-269] ^ d[511-266] ^ d[511-265] ^ d[511-261] ^ d[511-259] ^ d[511-257] ^ d[511-256] ^ d[511-255] ^ d[511-253] ^ d[511-251] ^ d[511-248] ^ d[511-246] ^ d[511-245] ^ d[511-244] ^ d[511-243] ^ d[511-242] ^ d[511-241] ^ d[511-235] ^ d[511-234] ^ d[511-230] ^ d[511-229] ^ d[511-228] ^ d[511-227] ^ d[511-222] ^ d[511-220] ^ d[511-219] ^ d[511-218] ^ d[511-217] ^ d[511-216] ^ d[511-215] ^ d[511-214] ^ d[511-210] ^ d[511-207] ^ d[511-206] ^ d[511-204] ^ d[511-201] ^ d[511-199] ^ d[511-197] ^ d[511-196] ^ d[511-194] ^ d[511-193] ^ d[511-192] ^ d[511-190] ^ d[511-188] ^ d[511-187] ^ d[511-185] ^ d[511-184] ^ d[511-181] ^ d[511-180] ^ d[511-177] ^ d[511-175] ^ d[511-170] ^ d[511-169] ^ d[511-168] ^ d[511-167] ^ d[511-165] ^ d[511-162] ^ d[511-158] ^ d[511-157] ^ d[511-156] ^ d[511-154] ^ d[511-153] ^ d[511-149] ^ d[511-145] ^ d[511-141] ^ d[511-137] ^ d[511-136] ^ d[511-134] ^ d[511-133] ^ d[511-128] ^ d[511-127] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-117] ^ d[511-116] ^ d[511-113] ^ d[511-111] ^ d[511-110] ^ d[511-109] ^ d[511-108] ^ d[511-105] ^ d[511-102] ^ d[511-101] ^ d[511-98] ^ d[511-97] ^ d[511-96] ^ d[511-94] ^ d[511-92] ^ d[511-91] ^ d[511-87] ^ d[511-86] ^ d[511-85] ^ d[511-82] ^ d[511-81] ^ d[511-77] ^ d[511-75] ^ d[511-74] ^ d[511-73] ^ d[511-71] ^ d[511-69] ^ d[511-68] ^ d[511-63] ^ d[511-61] ^ d[511-59] ^ d[511-57] ^ d[511-56] ^ d[511-54] ^ d[511-53] ^ d[511-52] ^ d[511-51] ^ d[511-50] ^ d[511-49] ^ d[511-47] ^ d[511-46] ^ d[511-42] ^ d[511-41] ^ d[511-31] ^ d[511-30] ^ d[511-27] ^ d[511-24] ^ d[511-21] ^ d[511-18] ^ d[511-17] ^ d[511-15] ^ d[511-13] ^ d[511-12] ^ d[511-9] ^ d[511-6] ^ d[511-5] ^ d[511-4] ^ d[511-2] ^ d[511-1] ^ d[511-0] ^ c[31-4] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-12] ^ c[31-13] ^ c[31-15] ^ c[31-16] ^ c[31-20] ^ c[31-21] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-30];
                stage_crc512_crc[18] <= d[511-511] ^ d[511-509] ^ d[511-508] ^ d[511-507] ^ d[511-506] ^ d[511-505] ^ d[511-502] ^ d[511-501] ^ d[511-497] ^ d[511-496] ^ d[511-494] ^ d[511-493] ^ d[511-489] ^ d[511-488] ^ d[511-487] ^ d[511-485] ^ d[511-478] ^ d[511-477] ^ d[511-474] ^ d[511-473] ^ d[511-472] ^ d[511-471] ^ d[511-467] ^ d[511-465] ^ d[511-463] ^ d[511-462] ^ d[511-461] ^ d[511-459] ^ d[511-458] ^ d[511-456] ^ d[511-454] ^ d[511-452] ^ d[511-451] ^ d[511-447] ^ d[511-445] ^ d[511-438] ^ d[511-437] ^ d[511-436] ^ d[511-431] ^ d[511-429] ^ d[511-428] ^ d[511-426] ^ d[511-424] ^ d[511-420] ^ d[511-419] ^ d[511-418] ^ d[511-417] ^ d[511-416] ^ d[511-415] ^ d[511-412] ^ d[511-410] ^ d[511-408] ^ d[511-407] ^ d[511-406] ^ d[511-403] ^ d[511-397] ^ d[511-396] ^ d[511-395] ^ d[511-392] ^ d[511-388] ^ d[511-387] ^ d[511-386] ^ d[511-385] ^ d[511-381] ^ d[511-380] ^ d[511-379] ^ d[511-376] ^ d[511-373] ^ d[511-371] ^ d[511-369] ^ d[511-368] ^ d[511-365] ^ d[511-364] ^ d[511-363] ^ d[511-361] ^ d[511-359] ^ d[511-358] ^ d[511-356] ^ d[511-355] ^ d[511-352] ^ d[511-342] ^ d[511-341] ^ d[511-340] ^ d[511-337] ^ d[511-336] ^ d[511-333] ^ d[511-331] ^ d[511-330] ^ d[511-327] ^ d[511-326] ^ d[511-325] ^ d[511-321] ^ d[511-319] ^ d[511-315] ^ d[511-314] ^ d[511-313] ^ d[511-312] ^ d[511-309] ^ d[511-307] ^ d[511-306] ^ d[511-304] ^ d[511-298] ^ d[511-292] ^ d[511-291] ^ d[511-281] ^ d[511-280] ^ d[511-279] ^ d[511-278] ^ d[511-276] ^ d[511-274] ^ d[511-270] ^ d[511-267] ^ d[511-266] ^ d[511-262] ^ d[511-260] ^ d[511-258] ^ d[511-257] ^ d[511-256] ^ d[511-254] ^ d[511-252] ^ d[511-249] ^ d[511-247] ^ d[511-246] ^ d[511-245] ^ d[511-244] ^ d[511-243] ^ d[511-242] ^ d[511-236] ^ d[511-235] ^ d[511-231] ^ d[511-230] ^ d[511-229] ^ d[511-228] ^ d[511-223] ^ d[511-221] ^ d[511-220] ^ d[511-219] ^ d[511-218] ^ d[511-217] ^ d[511-216] ^ d[511-215] ^ d[511-211] ^ d[511-208] ^ d[511-207] ^ d[511-205] ^ d[511-202] ^ d[511-200] ^ d[511-198] ^ d[511-197] ^ d[511-195] ^ d[511-194] ^ d[511-193] ^ d[511-191] ^ d[511-189] ^ d[511-188] ^ d[511-186] ^ d[511-185] ^ d[511-182] ^ d[511-181] ^ d[511-178] ^ d[511-176] ^ d[511-171] ^ d[511-170] ^ d[511-169] ^ d[511-168] ^ d[511-166] ^ d[511-163] ^ d[511-159] ^ d[511-158] ^ d[511-157] ^ d[511-155] ^ d[511-154] ^ d[511-150] ^ d[511-146] ^ d[511-142] ^ d[511-138] ^ d[511-137] ^ d[511-135] ^ d[511-134] ^ d[511-129] ^ d[511-128] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-118] ^ d[511-117] ^ d[511-114] ^ d[511-112] ^ d[511-111] ^ d[511-110] ^ d[511-109] ^ d[511-106] ^ d[511-103] ^ d[511-102] ^ d[511-99] ^ d[511-98] ^ d[511-97] ^ d[511-95] ^ d[511-93] ^ d[511-92] ^ d[511-88] ^ d[511-87] ^ d[511-86] ^ d[511-83] ^ d[511-82] ^ d[511-78] ^ d[511-76] ^ d[511-75] ^ d[511-74] ^ d[511-72] ^ d[511-70] ^ d[511-69] ^ d[511-64] ^ d[511-62] ^ d[511-60] ^ d[511-58] ^ d[511-57] ^ d[511-55] ^ d[511-54] ^ d[511-53] ^ d[511-52] ^ d[511-51] ^ d[511-50] ^ d[511-48] ^ d[511-47] ^ d[511-43] ^ d[511-42] ^ d[511-32] ^ d[511-31] ^ d[511-28] ^ d[511-25] ^ d[511-22] ^ d[511-19] ^ d[511-18] ^ d[511-16] ^ d[511-14] ^ d[511-13] ^ d[511-10] ^ d[511-7] ^ d[511-6] ^ d[511-5] ^ d[511-3] ^ d[511-2] ^ d[511-1] ^ c[31-5] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-13] ^ c[31-14] ^ c[31-16] ^ c[31-17] ^ c[31-21] ^ c[31-22] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-31];
                stage_crc512_crc[17] <= d[511-510] ^ d[511-509] ^ d[511-508] ^ d[511-507] ^ d[511-506] ^ d[511-503] ^ d[511-502] ^ d[511-498] ^ d[511-497] ^ d[511-495] ^ d[511-494] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-486] ^ d[511-479] ^ d[511-478] ^ d[511-475] ^ d[511-474] ^ d[511-473] ^ d[511-472] ^ d[511-468] ^ d[511-466] ^ d[511-464] ^ d[511-463] ^ d[511-462] ^ d[511-460] ^ d[511-459] ^ d[511-457] ^ d[511-455] ^ d[511-453] ^ d[511-452] ^ d[511-448] ^ d[511-446] ^ d[511-439] ^ d[511-438] ^ d[511-437] ^ d[511-432] ^ d[511-430] ^ d[511-429] ^ d[511-427] ^ d[511-425] ^ d[511-421] ^ d[511-420] ^ d[511-419] ^ d[511-418] ^ d[511-417] ^ d[511-416] ^ d[511-413] ^ d[511-411] ^ d[511-409] ^ d[511-408] ^ d[511-407] ^ d[511-404] ^ d[511-398] ^ d[511-397] ^ d[511-396] ^ d[511-393] ^ d[511-389] ^ d[511-388] ^ d[511-387] ^ d[511-386] ^ d[511-382] ^ d[511-381] ^ d[511-380] ^ d[511-377] ^ d[511-374] ^ d[511-372] ^ d[511-370] ^ d[511-369] ^ d[511-366] ^ d[511-365] ^ d[511-364] ^ d[511-362] ^ d[511-360] ^ d[511-359] ^ d[511-357] ^ d[511-356] ^ d[511-353] ^ d[511-343] ^ d[511-342] ^ d[511-341] ^ d[511-338] ^ d[511-337] ^ d[511-334] ^ d[511-332] ^ d[511-331] ^ d[511-328] ^ d[511-327] ^ d[511-326] ^ d[511-322] ^ d[511-320] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-313] ^ d[511-310] ^ d[511-308] ^ d[511-307] ^ d[511-305] ^ d[511-299] ^ d[511-293] ^ d[511-292] ^ d[511-282] ^ d[511-281] ^ d[511-280] ^ d[511-279] ^ d[511-277] ^ d[511-275] ^ d[511-271] ^ d[511-268] ^ d[511-267] ^ d[511-263] ^ d[511-261] ^ d[511-259] ^ d[511-258] ^ d[511-257] ^ d[511-255] ^ d[511-253] ^ d[511-250] ^ d[511-248] ^ d[511-247] ^ d[511-246] ^ d[511-245] ^ d[511-244] ^ d[511-243] ^ d[511-237] ^ d[511-236] ^ d[511-232] ^ d[511-231] ^ d[511-230] ^ d[511-229] ^ d[511-224] ^ d[511-222] ^ d[511-221] ^ d[511-220] ^ d[511-219] ^ d[511-218] ^ d[511-217] ^ d[511-216] ^ d[511-212] ^ d[511-209] ^ d[511-208] ^ d[511-206] ^ d[511-203] ^ d[511-201] ^ d[511-199] ^ d[511-198] ^ d[511-196] ^ d[511-195] ^ d[511-194] ^ d[511-192] ^ d[511-190] ^ d[511-189] ^ d[511-187] ^ d[511-186] ^ d[511-183] ^ d[511-182] ^ d[511-179] ^ d[511-177] ^ d[511-172] ^ d[511-171] ^ d[511-170] ^ d[511-169] ^ d[511-167] ^ d[511-164] ^ d[511-160] ^ d[511-159] ^ d[511-158] ^ d[511-156] ^ d[511-155] ^ d[511-151] ^ d[511-147] ^ d[511-143] ^ d[511-139] ^ d[511-138] ^ d[511-136] ^ d[511-135] ^ d[511-130] ^ d[511-129] ^ d[511-124] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-119] ^ d[511-118] ^ d[511-115] ^ d[511-113] ^ d[511-112] ^ d[511-111] ^ d[511-110] ^ d[511-107] ^ d[511-104] ^ d[511-103] ^ d[511-100] ^ d[511-99] ^ d[511-98] ^ d[511-96] ^ d[511-94] ^ d[511-93] ^ d[511-89] ^ d[511-88] ^ d[511-87] ^ d[511-84] ^ d[511-83] ^ d[511-79] ^ d[511-77] ^ d[511-76] ^ d[511-75] ^ d[511-73] ^ d[511-71] ^ d[511-70] ^ d[511-65] ^ d[511-63] ^ d[511-61] ^ d[511-59] ^ d[511-58] ^ d[511-56] ^ d[511-55] ^ d[511-54] ^ d[511-53] ^ d[511-52] ^ d[511-51] ^ d[511-49] ^ d[511-48] ^ d[511-44] ^ d[511-43] ^ d[511-33] ^ d[511-32] ^ d[511-29] ^ d[511-26] ^ d[511-23] ^ d[511-20] ^ d[511-19] ^ d[511-17] ^ d[511-15] ^ d[511-14] ^ d[511-11] ^ d[511-8] ^ d[511-7] ^ d[511-6] ^ d[511-4] ^ d[511-3] ^ d[511-2] ^ c[31-6] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-14] ^ c[31-15] ^ c[31-17] ^ c[31-18] ^ c[31-22] ^ c[31-23] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30];
                stage_crc512_crc[16] <= d[511-511] ^ d[511-510] ^ d[511-509] ^ d[511-508] ^ d[511-507] ^ d[511-504] ^ d[511-503] ^ d[511-499] ^ d[511-498] ^ d[511-496] ^ d[511-495] ^ d[511-491] ^ d[511-490] ^ d[511-489] ^ d[511-487] ^ d[511-480] ^ d[511-479] ^ d[511-476] ^ d[511-475] ^ d[511-474] ^ d[511-473] ^ d[511-469] ^ d[511-467] ^ d[511-465] ^ d[511-464] ^ d[511-463] ^ d[511-461] ^ d[511-460] ^ d[511-458] ^ d[511-456] ^ d[511-454] ^ d[511-453] ^ d[511-449] ^ d[511-447] ^ d[511-440] ^ d[511-439] ^ d[511-438] ^ d[511-433] ^ d[511-431] ^ d[511-430] ^ d[511-428] ^ d[511-426] ^ d[511-422] ^ d[511-421] ^ d[511-420] ^ d[511-419] ^ d[511-418] ^ d[511-417] ^ d[511-414] ^ d[511-412] ^ d[511-410] ^ d[511-409] ^ d[511-408] ^ d[511-405] ^ d[511-399] ^ d[511-398] ^ d[511-397] ^ d[511-394] ^ d[511-390] ^ d[511-389] ^ d[511-388] ^ d[511-387] ^ d[511-383] ^ d[511-382] ^ d[511-381] ^ d[511-378] ^ d[511-375] ^ d[511-373] ^ d[511-371] ^ d[511-370] ^ d[511-367] ^ d[511-366] ^ d[511-365] ^ d[511-363] ^ d[511-361] ^ d[511-360] ^ d[511-358] ^ d[511-357] ^ d[511-354] ^ d[511-344] ^ d[511-343] ^ d[511-342] ^ d[511-339] ^ d[511-338] ^ d[511-335] ^ d[511-333] ^ d[511-332] ^ d[511-329] ^ d[511-328] ^ d[511-327] ^ d[511-323] ^ d[511-321] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-311] ^ d[511-309] ^ d[511-308] ^ d[511-306] ^ d[511-300] ^ d[511-294] ^ d[511-293] ^ d[511-283] ^ d[511-282] ^ d[511-281] ^ d[511-280] ^ d[511-278] ^ d[511-276] ^ d[511-272] ^ d[511-269] ^ d[511-268] ^ d[511-264] ^ d[511-262] ^ d[511-260] ^ d[511-259] ^ d[511-258] ^ d[511-256] ^ d[511-254] ^ d[511-251] ^ d[511-249] ^ d[511-248] ^ d[511-247] ^ d[511-246] ^ d[511-245] ^ d[511-244] ^ d[511-238] ^ d[511-237] ^ d[511-233] ^ d[511-232] ^ d[511-231] ^ d[511-230] ^ d[511-225] ^ d[511-223] ^ d[511-222] ^ d[511-221] ^ d[511-220] ^ d[511-219] ^ d[511-218] ^ d[511-217] ^ d[511-213] ^ d[511-210] ^ d[511-209] ^ d[511-207] ^ d[511-204] ^ d[511-202] ^ d[511-200] ^ d[511-199] ^ d[511-197] ^ d[511-196] ^ d[511-195] ^ d[511-193] ^ d[511-191] ^ d[511-190] ^ d[511-188] ^ d[511-187] ^ d[511-184] ^ d[511-183] ^ d[511-180] ^ d[511-178] ^ d[511-173] ^ d[511-172] ^ d[511-171] ^ d[511-170] ^ d[511-168] ^ d[511-165] ^ d[511-161] ^ d[511-160] ^ d[511-159] ^ d[511-157] ^ d[511-156] ^ d[511-152] ^ d[511-148] ^ d[511-144] ^ d[511-140] ^ d[511-139] ^ d[511-137] ^ d[511-136] ^ d[511-131] ^ d[511-130] ^ d[511-125] ^ d[511-124] ^ d[511-123] ^ d[511-122] ^ d[511-120] ^ d[511-119] ^ d[511-116] ^ d[511-114] ^ d[511-113] ^ d[511-112] ^ d[511-111] ^ d[511-108] ^ d[511-105] ^ d[511-104] ^ d[511-101] ^ d[511-100] ^ d[511-99] ^ d[511-97] ^ d[511-95] ^ d[511-94] ^ d[511-90] ^ d[511-89] ^ d[511-88] ^ d[511-85] ^ d[511-84] ^ d[511-80] ^ d[511-78] ^ d[511-77] ^ d[511-76] ^ d[511-74] ^ d[511-72] ^ d[511-71] ^ d[511-66] ^ d[511-64] ^ d[511-62] ^ d[511-60] ^ d[511-59] ^ d[511-57] ^ d[511-56] ^ d[511-55] ^ d[511-54] ^ d[511-53] ^ d[511-52] ^ d[511-50] ^ d[511-49] ^ d[511-45] ^ d[511-44] ^ d[511-34] ^ d[511-33] ^ d[511-30] ^ d[511-27] ^ d[511-24] ^ d[511-21] ^ d[511-20] ^ d[511-18] ^ d[511-16] ^ d[511-15] ^ d[511-12] ^ d[511-9] ^ d[511-8] ^ d[511-7] ^ d[511-5] ^ d[511-4] ^ d[511-3] ^ c[31-0] ^ c[31-7] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-15] ^ c[31-16] ^ c[31-18] ^ c[31-19] ^ c[31-23] ^ c[31-24] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc512_crc[15] <= d[511-509] ^ d[511-507] ^ d[511-506] ^ d[511-505] ^ d[511-504] ^ d[511-502] ^ d[511-501] ^ d[511-499] ^ d[511-497] ^ d[511-496] ^ d[511-495] ^ d[511-494] ^ d[511-493] ^ d[511-489] ^ d[511-486] ^ d[511-483] ^ d[511-482] ^ d[511-479] ^ d[511-475] ^ d[511-474] ^ d[511-472] ^ d[511-466] ^ d[511-459] ^ d[511-458] ^ d[511-457] ^ d[511-455] ^ d[511-454] ^ d[511-452] ^ d[511-449] ^ d[511-444] ^ d[511-441] ^ d[511-440] ^ d[511-439] ^ d[511-437] ^ d[511-436] ^ d[511-433] ^ d[511-432] ^ d[511-431] ^ d[511-429] ^ d[511-427] ^ d[511-424] ^ d[511-423] ^ d[511-421] ^ d[511-420] ^ d[511-416] ^ d[511-415] ^ d[511-414] ^ d[511-413] ^ d[511-412] ^ d[511-411] ^ d[511-410] ^ d[511-408] ^ d[511-407] ^ d[511-406] ^ d[511-405] ^ d[511-404] ^ d[511-396] ^ d[511-395] ^ d[511-393] ^ d[511-392] ^ d[511-389] ^ d[511-387] ^ d[511-386] ^ d[511-384] ^ d[511-383] ^ d[511-382] ^ d[511-381] ^ d[511-379] ^ d[511-378] ^ d[511-371] ^ d[511-369] ^ d[511-367] ^ d[511-364] ^ d[511-363] ^ d[511-361] ^ d[511-357] ^ d[511-355] ^ d[511-353] ^ d[511-349] ^ d[511-348] ^ d[511-347] ^ d[511-343] ^ d[511-342] ^ d[511-341] ^ d[511-340] ^ d[511-338] ^ d[511-337] ^ d[511-336] ^ d[511-335] ^ d[511-330] ^ d[511-329] ^ d[511-327] ^ d[511-324] ^ d[511-321] ^ d[511-320] ^ d[511-319] ^ d[511-316] ^ d[511-307] ^ d[511-305] ^ d[511-303] ^ d[511-302] ^ d[511-301] ^ d[511-300] ^ d[511-299] ^ d[511-298] ^ d[511-297] ^ d[511-296] ^ d[511-292] ^ d[511-290] ^ d[511-288] ^ d[511-287] ^ d[511-286] ^ d[511-284] ^ d[511-282] ^ d[511-281] ^ d[511-276] ^ d[511-274] ^ d[511-270] ^ d[511-268] ^ d[511-264] ^ d[511-263] ^ d[511-260] ^ d[511-250] ^ d[511-249] ^ d[511-247] ^ d[511-246] ^ d[511-245] ^ d[511-243] ^ d[511-239] ^ d[511-238] ^ d[511-237] ^ d[511-233] ^ d[511-232] ^ d[511-231] ^ d[511-230] ^ d[511-228] ^ d[511-227] ^ d[511-223] ^ d[511-222] ^ d[511-221] ^ d[511-220] ^ d[511-219] ^ d[511-218] ^ d[511-216] ^ d[511-212] ^ d[511-211] ^ d[511-209] ^ d[511-207] ^ d[511-205] ^ d[511-202] ^ d[511-200] ^ d[511-199] ^ d[511-196] ^ d[511-193] ^ d[511-190] ^ d[511-189] ^ d[511-186] ^ d[511-185] ^ d[511-184] ^ d[511-183] ^ d[511-182] ^ d[511-181] ^ d[511-179] ^ d[511-174] ^ d[511-173] ^ d[511-170] ^ d[511-167] ^ d[511-160] ^ d[511-157] ^ d[511-156] ^ d[511-155] ^ d[511-153] ^ d[511-151] ^ d[511-145] ^ d[511-144] ^ d[511-143] ^ d[511-141] ^ d[511-140] ^ d[511-138] ^ d[511-136] ^ d[511-135] ^ d[511-134] ^ d[511-131] ^ d[511-128] ^ d[511-127] ^ d[511-124] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-118] ^ d[511-116] ^ d[511-115] ^ d[511-112] ^ d[511-111] ^ d[511-110] ^ d[511-109] ^ d[511-105] ^ d[511-104] ^ d[511-103] ^ d[511-102] ^ d[511-100] ^ d[511-99] ^ d[511-97] ^ d[511-94] ^ d[511-91] ^ d[511-90] ^ d[511-89] ^ d[511-87] ^ d[511-86] ^ d[511-84] ^ d[511-83] ^ d[511-82] ^ d[511-78] ^ d[511-77] ^ d[511-75] ^ d[511-68] ^ d[511-66] ^ d[511-57] ^ d[511-56] ^ d[511-51] ^ d[511-48] ^ d[511-47] ^ d[511-46] ^ d[511-44] ^ d[511-37] ^ d[511-35] ^ d[511-32] ^ d[511-30] ^ d[511-29] ^ d[511-26] ^ d[511-24] ^ d[511-22] ^ d[511-21] ^ d[511-19] ^ d[511-17] ^ d[511-13] ^ d[511-12] ^ d[511-8] ^ d[511-5] ^ d[511-4] ^ d[511-0] ^ c[31-2] ^ c[31-3] ^ c[31-6] ^ c[31-9] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-19] ^ c[31-21] ^ c[31-22] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-29];
                stage_crc512_crc[14] <= d[511-510] ^ d[511-508] ^ d[511-507] ^ d[511-506] ^ d[511-505] ^ d[511-503] ^ d[511-502] ^ d[511-500] ^ d[511-498] ^ d[511-497] ^ d[511-496] ^ d[511-495] ^ d[511-494] ^ d[511-490] ^ d[511-487] ^ d[511-484] ^ d[511-483] ^ d[511-480] ^ d[511-476] ^ d[511-475] ^ d[511-473] ^ d[511-467] ^ d[511-460] ^ d[511-459] ^ d[511-458] ^ d[511-456] ^ d[511-455] ^ d[511-453] ^ d[511-450] ^ d[511-445] ^ d[511-442] ^ d[511-441] ^ d[511-440] ^ d[511-438] ^ d[511-437] ^ d[511-434] ^ d[511-433] ^ d[511-432] ^ d[511-430] ^ d[511-428] ^ d[511-425] ^ d[511-424] ^ d[511-422] ^ d[511-421] ^ d[511-417] ^ d[511-416] ^ d[511-415] ^ d[511-414] ^ d[511-413] ^ d[511-412] ^ d[511-411] ^ d[511-409] ^ d[511-408] ^ d[511-407] ^ d[511-406] ^ d[511-405] ^ d[511-397] ^ d[511-396] ^ d[511-394] ^ d[511-393] ^ d[511-390] ^ d[511-388] ^ d[511-387] ^ d[511-385] ^ d[511-384] ^ d[511-383] ^ d[511-382] ^ d[511-380] ^ d[511-379] ^ d[511-372] ^ d[511-370] ^ d[511-368] ^ d[511-365] ^ d[511-364] ^ d[511-362] ^ d[511-358] ^ d[511-356] ^ d[511-354] ^ d[511-350] ^ d[511-349] ^ d[511-348] ^ d[511-344] ^ d[511-343] ^ d[511-342] ^ d[511-341] ^ d[511-339] ^ d[511-338] ^ d[511-337] ^ d[511-336] ^ d[511-331] ^ d[511-330] ^ d[511-328] ^ d[511-325] ^ d[511-322] ^ d[511-321] ^ d[511-320] ^ d[511-317] ^ d[511-308] ^ d[511-306] ^ d[511-304] ^ d[511-303] ^ d[511-302] ^ d[511-301] ^ d[511-300] ^ d[511-299] ^ d[511-298] ^ d[511-297] ^ d[511-293] ^ d[511-291] ^ d[511-289] ^ d[511-288] ^ d[511-287] ^ d[511-285] ^ d[511-283] ^ d[511-282] ^ d[511-277] ^ d[511-275] ^ d[511-271] ^ d[511-269] ^ d[511-265] ^ d[511-264] ^ d[511-261] ^ d[511-251] ^ d[511-250] ^ d[511-248] ^ d[511-247] ^ d[511-246] ^ d[511-244] ^ d[511-240] ^ d[511-239] ^ d[511-238] ^ d[511-234] ^ d[511-233] ^ d[511-232] ^ d[511-231] ^ d[511-229] ^ d[511-228] ^ d[511-224] ^ d[511-223] ^ d[511-222] ^ d[511-221] ^ d[511-220] ^ d[511-219] ^ d[511-217] ^ d[511-213] ^ d[511-212] ^ d[511-210] ^ d[511-208] ^ d[511-206] ^ d[511-203] ^ d[511-201] ^ d[511-200] ^ d[511-197] ^ d[511-194] ^ d[511-191] ^ d[511-190] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-184] ^ d[511-183] ^ d[511-182] ^ d[511-180] ^ d[511-175] ^ d[511-174] ^ d[511-171] ^ d[511-168] ^ d[511-161] ^ d[511-158] ^ d[511-157] ^ d[511-156] ^ d[511-154] ^ d[511-152] ^ d[511-146] ^ d[511-145] ^ d[511-144] ^ d[511-142] ^ d[511-141] ^ d[511-139] ^ d[511-137] ^ d[511-136] ^ d[511-135] ^ d[511-132] ^ d[511-129] ^ d[511-128] ^ d[511-125] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-117] ^ d[511-116] ^ d[511-113] ^ d[511-112] ^ d[511-111] ^ d[511-110] ^ d[511-106] ^ d[511-105] ^ d[511-104] ^ d[511-103] ^ d[511-101] ^ d[511-100] ^ d[511-98] ^ d[511-95] ^ d[511-92] ^ d[511-91] ^ d[511-90] ^ d[511-88] ^ d[511-87] ^ d[511-85] ^ d[511-84] ^ d[511-83] ^ d[511-79] ^ d[511-78] ^ d[511-76] ^ d[511-69] ^ d[511-67] ^ d[511-58] ^ d[511-57] ^ d[511-52] ^ d[511-49] ^ d[511-48] ^ d[511-47] ^ d[511-45] ^ d[511-38] ^ d[511-36] ^ d[511-33] ^ d[511-31] ^ d[511-30] ^ d[511-27] ^ d[511-25] ^ d[511-23] ^ d[511-22] ^ d[511-20] ^ d[511-18] ^ d[511-14] ^ d[511-13] ^ d[511-9] ^ d[511-6] ^ d[511-5] ^ d[511-1] ^ c[31-0] ^ c[31-3] ^ c[31-4] ^ c[31-7] ^ c[31-10] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-20] ^ c[31-22] ^ c[31-23] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-30];
                stage_crc512_crc[13] <= d[511-511] ^ d[511-509] ^ d[511-508] ^ d[511-507] ^ d[511-506] ^ d[511-504] ^ d[511-503] ^ d[511-501] ^ d[511-499] ^ d[511-498] ^ d[511-497] ^ d[511-496] ^ d[511-495] ^ d[511-491] ^ d[511-488] ^ d[511-485] ^ d[511-484] ^ d[511-481] ^ d[511-477] ^ d[511-476] ^ d[511-474] ^ d[511-468] ^ d[511-461] ^ d[511-460] ^ d[511-459] ^ d[511-457] ^ d[511-456] ^ d[511-454] ^ d[511-451] ^ d[511-446] ^ d[511-443] ^ d[511-442] ^ d[511-441] ^ d[511-439] ^ d[511-438] ^ d[511-435] ^ d[511-434] ^ d[511-433] ^ d[511-431] ^ d[511-429] ^ d[511-426] ^ d[511-425] ^ d[511-423] ^ d[511-422] ^ d[511-418] ^ d[511-417] ^ d[511-416] ^ d[511-415] ^ d[511-414] ^ d[511-413] ^ d[511-412] ^ d[511-410] ^ d[511-409] ^ d[511-408] ^ d[511-407] ^ d[511-406] ^ d[511-398] ^ d[511-397] ^ d[511-395] ^ d[511-394] ^ d[511-391] ^ d[511-389] ^ d[511-388] ^ d[511-386] ^ d[511-385] ^ d[511-384] ^ d[511-383] ^ d[511-381] ^ d[511-380] ^ d[511-373] ^ d[511-371] ^ d[511-369] ^ d[511-366] ^ d[511-365] ^ d[511-363] ^ d[511-359] ^ d[511-357] ^ d[511-355] ^ d[511-351] ^ d[511-350] ^ d[511-349] ^ d[511-345] ^ d[511-344] ^ d[511-343] ^ d[511-342] ^ d[511-340] ^ d[511-339] ^ d[511-338] ^ d[511-337] ^ d[511-332] ^ d[511-331] ^ d[511-329] ^ d[511-326] ^ d[511-323] ^ d[511-322] ^ d[511-321] ^ d[511-318] ^ d[511-309] ^ d[511-307] ^ d[511-305] ^ d[511-304] ^ d[511-303] ^ d[511-302] ^ d[511-301] ^ d[511-300] ^ d[511-299] ^ d[511-298] ^ d[511-294] ^ d[511-292] ^ d[511-290] ^ d[511-289] ^ d[511-288] ^ d[511-286] ^ d[511-284] ^ d[511-283] ^ d[511-278] ^ d[511-276] ^ d[511-272] ^ d[511-270] ^ d[511-266] ^ d[511-265] ^ d[511-262] ^ d[511-252] ^ d[511-251] ^ d[511-249] ^ d[511-248] ^ d[511-247] ^ d[511-245] ^ d[511-241] ^ d[511-240] ^ d[511-239] ^ d[511-235] ^ d[511-234] ^ d[511-233] ^ d[511-232] ^ d[511-230] ^ d[511-229] ^ d[511-225] ^ d[511-224] ^ d[511-223] ^ d[511-222] ^ d[511-221] ^ d[511-220] ^ d[511-218] ^ d[511-214] ^ d[511-213] ^ d[511-211] ^ d[511-209] ^ d[511-207] ^ d[511-204] ^ d[511-202] ^ d[511-201] ^ d[511-198] ^ d[511-195] ^ d[511-192] ^ d[511-191] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-184] ^ d[511-183] ^ d[511-181] ^ d[511-176] ^ d[511-175] ^ d[511-172] ^ d[511-169] ^ d[511-162] ^ d[511-159] ^ d[511-158] ^ d[511-157] ^ d[511-155] ^ d[511-153] ^ d[511-147] ^ d[511-146] ^ d[511-145] ^ d[511-143] ^ d[511-142] ^ d[511-140] ^ d[511-138] ^ d[511-137] ^ d[511-136] ^ d[511-133] ^ d[511-130] ^ d[511-129] ^ d[511-126] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-118] ^ d[511-117] ^ d[511-114] ^ d[511-113] ^ d[511-112] ^ d[511-111] ^ d[511-107] ^ d[511-106] ^ d[511-105] ^ d[511-104] ^ d[511-102] ^ d[511-101] ^ d[511-99] ^ d[511-96] ^ d[511-93] ^ d[511-92] ^ d[511-91] ^ d[511-89] ^ d[511-88] ^ d[511-86] ^ d[511-85] ^ d[511-84] ^ d[511-80] ^ d[511-79] ^ d[511-77] ^ d[511-70] ^ d[511-68] ^ d[511-59] ^ d[511-58] ^ d[511-53] ^ d[511-50] ^ d[511-49] ^ d[511-48] ^ d[511-46] ^ d[511-39] ^ d[511-37] ^ d[511-34] ^ d[511-32] ^ d[511-31] ^ d[511-28] ^ d[511-26] ^ d[511-24] ^ d[511-23] ^ d[511-21] ^ d[511-19] ^ d[511-15] ^ d[511-14] ^ d[511-10] ^ d[511-7] ^ d[511-6] ^ d[511-2] ^ c[31-1] ^ c[31-4] ^ c[31-5] ^ c[31-8] ^ c[31-11] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-19] ^ c[31-21] ^ c[31-23] ^ c[31-24] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-31];
                stage_crc512_crc[12] <= d[511-510] ^ d[511-509] ^ d[511-508] ^ d[511-507] ^ d[511-505] ^ d[511-504] ^ d[511-502] ^ d[511-500] ^ d[511-499] ^ d[511-498] ^ d[511-497] ^ d[511-496] ^ d[511-492] ^ d[511-489] ^ d[511-486] ^ d[511-485] ^ d[511-482] ^ d[511-478] ^ d[511-477] ^ d[511-475] ^ d[511-469] ^ d[511-462] ^ d[511-461] ^ d[511-460] ^ d[511-458] ^ d[511-457] ^ d[511-455] ^ d[511-452] ^ d[511-447] ^ d[511-444] ^ d[511-443] ^ d[511-442] ^ d[511-440] ^ d[511-439] ^ d[511-436] ^ d[511-435] ^ d[511-434] ^ d[511-432] ^ d[511-430] ^ d[511-427] ^ d[511-426] ^ d[511-424] ^ d[511-423] ^ d[511-419] ^ d[511-418] ^ d[511-417] ^ d[511-416] ^ d[511-415] ^ d[511-414] ^ d[511-413] ^ d[511-411] ^ d[511-410] ^ d[511-409] ^ d[511-408] ^ d[511-407] ^ d[511-399] ^ d[511-398] ^ d[511-396] ^ d[511-395] ^ d[511-392] ^ d[511-390] ^ d[511-389] ^ d[511-387] ^ d[511-386] ^ d[511-385] ^ d[511-384] ^ d[511-382] ^ d[511-381] ^ d[511-374] ^ d[511-372] ^ d[511-370] ^ d[511-367] ^ d[511-366] ^ d[511-364] ^ d[511-360] ^ d[511-358] ^ d[511-356] ^ d[511-352] ^ d[511-351] ^ d[511-350] ^ d[511-346] ^ d[511-345] ^ d[511-344] ^ d[511-343] ^ d[511-341] ^ d[511-340] ^ d[511-339] ^ d[511-338] ^ d[511-333] ^ d[511-332] ^ d[511-330] ^ d[511-327] ^ d[511-324] ^ d[511-323] ^ d[511-322] ^ d[511-319] ^ d[511-310] ^ d[511-308] ^ d[511-306] ^ d[511-305] ^ d[511-304] ^ d[511-303] ^ d[511-302] ^ d[511-301] ^ d[511-300] ^ d[511-299] ^ d[511-295] ^ d[511-293] ^ d[511-291] ^ d[511-290] ^ d[511-289] ^ d[511-287] ^ d[511-285] ^ d[511-284] ^ d[511-279] ^ d[511-277] ^ d[511-273] ^ d[511-271] ^ d[511-267] ^ d[511-266] ^ d[511-263] ^ d[511-253] ^ d[511-252] ^ d[511-250] ^ d[511-249] ^ d[511-248] ^ d[511-246] ^ d[511-242] ^ d[511-241] ^ d[511-240] ^ d[511-236] ^ d[511-235] ^ d[511-234] ^ d[511-233] ^ d[511-231] ^ d[511-230] ^ d[511-226] ^ d[511-225] ^ d[511-224] ^ d[511-223] ^ d[511-222] ^ d[511-221] ^ d[511-219] ^ d[511-215] ^ d[511-214] ^ d[511-212] ^ d[511-210] ^ d[511-208] ^ d[511-205] ^ d[511-203] ^ d[511-202] ^ d[511-199] ^ d[511-196] ^ d[511-193] ^ d[511-192] ^ d[511-189] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-184] ^ d[511-182] ^ d[511-177] ^ d[511-176] ^ d[511-173] ^ d[511-170] ^ d[511-163] ^ d[511-160] ^ d[511-159] ^ d[511-158] ^ d[511-156] ^ d[511-154] ^ d[511-148] ^ d[511-147] ^ d[511-146] ^ d[511-144] ^ d[511-143] ^ d[511-141] ^ d[511-139] ^ d[511-138] ^ d[511-137] ^ d[511-134] ^ d[511-131] ^ d[511-130] ^ d[511-127] ^ d[511-124] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-119] ^ d[511-118] ^ d[511-115] ^ d[511-114] ^ d[511-113] ^ d[511-112] ^ d[511-108] ^ d[511-107] ^ d[511-106] ^ d[511-105] ^ d[511-103] ^ d[511-102] ^ d[511-100] ^ d[511-97] ^ d[511-94] ^ d[511-93] ^ d[511-92] ^ d[511-90] ^ d[511-89] ^ d[511-87] ^ d[511-86] ^ d[511-85] ^ d[511-81] ^ d[511-80] ^ d[511-78] ^ d[511-71] ^ d[511-69] ^ d[511-60] ^ d[511-59] ^ d[511-54] ^ d[511-51] ^ d[511-50] ^ d[511-49] ^ d[511-47] ^ d[511-40] ^ d[511-38] ^ d[511-35] ^ d[511-33] ^ d[511-32] ^ d[511-29] ^ d[511-27] ^ d[511-25] ^ d[511-24] ^ d[511-22] ^ d[511-20] ^ d[511-16] ^ d[511-15] ^ d[511-11] ^ d[511-8] ^ d[511-7] ^ d[511-3] ^ c[31-2] ^ c[31-5] ^ c[31-6] ^ c[31-9] ^ c[31-12] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-19] ^ c[31-20] ^ c[31-22] ^ c[31-24] ^ c[31-25] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30];
                stage_crc512_crc[11] <= d[511-511] ^ d[511-510] ^ d[511-509] ^ d[511-508] ^ d[511-506] ^ d[511-505] ^ d[511-503] ^ d[511-501] ^ d[511-500] ^ d[511-499] ^ d[511-498] ^ d[511-497] ^ d[511-493] ^ d[511-490] ^ d[511-487] ^ d[511-486] ^ d[511-483] ^ d[511-479] ^ d[511-478] ^ d[511-476] ^ d[511-470] ^ d[511-463] ^ d[511-462] ^ d[511-461] ^ d[511-459] ^ d[511-458] ^ d[511-456] ^ d[511-453] ^ d[511-448] ^ d[511-445] ^ d[511-444] ^ d[511-443] ^ d[511-441] ^ d[511-440] ^ d[511-437] ^ d[511-436] ^ d[511-435] ^ d[511-433] ^ d[511-431] ^ d[511-428] ^ d[511-427] ^ d[511-425] ^ d[511-424] ^ d[511-420] ^ d[511-419] ^ d[511-418] ^ d[511-417] ^ d[511-416] ^ d[511-415] ^ d[511-414] ^ d[511-412] ^ d[511-411] ^ d[511-410] ^ d[511-409] ^ d[511-408] ^ d[511-400] ^ d[511-399] ^ d[511-397] ^ d[511-396] ^ d[511-393] ^ d[511-391] ^ d[511-390] ^ d[511-388] ^ d[511-387] ^ d[511-386] ^ d[511-385] ^ d[511-383] ^ d[511-382] ^ d[511-375] ^ d[511-373] ^ d[511-371] ^ d[511-368] ^ d[511-367] ^ d[511-365] ^ d[511-361] ^ d[511-359] ^ d[511-357] ^ d[511-353] ^ d[511-352] ^ d[511-351] ^ d[511-347] ^ d[511-346] ^ d[511-345] ^ d[511-344] ^ d[511-342] ^ d[511-341] ^ d[511-340] ^ d[511-339] ^ d[511-334] ^ d[511-333] ^ d[511-331] ^ d[511-328] ^ d[511-325] ^ d[511-324] ^ d[511-323] ^ d[511-320] ^ d[511-311] ^ d[511-309] ^ d[511-307] ^ d[511-306] ^ d[511-305] ^ d[511-304] ^ d[511-303] ^ d[511-302] ^ d[511-301] ^ d[511-300] ^ d[511-296] ^ d[511-294] ^ d[511-292] ^ d[511-291] ^ d[511-290] ^ d[511-288] ^ d[511-286] ^ d[511-285] ^ d[511-280] ^ d[511-278] ^ d[511-274] ^ d[511-272] ^ d[511-268] ^ d[511-267] ^ d[511-264] ^ d[511-254] ^ d[511-253] ^ d[511-251] ^ d[511-250] ^ d[511-249] ^ d[511-247] ^ d[511-243] ^ d[511-242] ^ d[511-241] ^ d[511-237] ^ d[511-236] ^ d[511-235] ^ d[511-234] ^ d[511-232] ^ d[511-231] ^ d[511-227] ^ d[511-226] ^ d[511-225] ^ d[511-224] ^ d[511-223] ^ d[511-222] ^ d[511-220] ^ d[511-216] ^ d[511-215] ^ d[511-213] ^ d[511-211] ^ d[511-209] ^ d[511-206] ^ d[511-204] ^ d[511-203] ^ d[511-200] ^ d[511-197] ^ d[511-194] ^ d[511-193] ^ d[511-190] ^ d[511-189] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-183] ^ d[511-178] ^ d[511-177] ^ d[511-174] ^ d[511-171] ^ d[511-164] ^ d[511-161] ^ d[511-160] ^ d[511-159] ^ d[511-157] ^ d[511-155] ^ d[511-149] ^ d[511-148] ^ d[511-147] ^ d[511-145] ^ d[511-144] ^ d[511-142] ^ d[511-140] ^ d[511-139] ^ d[511-138] ^ d[511-135] ^ d[511-132] ^ d[511-131] ^ d[511-128] ^ d[511-125] ^ d[511-124] ^ d[511-123] ^ d[511-122] ^ d[511-120] ^ d[511-119] ^ d[511-116] ^ d[511-115] ^ d[511-114] ^ d[511-113] ^ d[511-109] ^ d[511-108] ^ d[511-107] ^ d[511-106] ^ d[511-104] ^ d[511-103] ^ d[511-101] ^ d[511-98] ^ d[511-95] ^ d[511-94] ^ d[511-93] ^ d[511-91] ^ d[511-90] ^ d[511-88] ^ d[511-87] ^ d[511-86] ^ d[511-82] ^ d[511-81] ^ d[511-79] ^ d[511-72] ^ d[511-70] ^ d[511-61] ^ d[511-60] ^ d[511-55] ^ d[511-52] ^ d[511-51] ^ d[511-50] ^ d[511-48] ^ d[511-41] ^ d[511-39] ^ d[511-36] ^ d[511-34] ^ d[511-33] ^ d[511-30] ^ d[511-28] ^ d[511-26] ^ d[511-25] ^ d[511-23] ^ d[511-21] ^ d[511-17] ^ d[511-16] ^ d[511-12] ^ d[511-9] ^ d[511-8] ^ d[511-4] ^ c[31-3] ^ c[31-6] ^ c[31-7] ^ c[31-10] ^ c[31-13] ^ c[31-17] ^ c[31-18] ^ c[31-19] ^ c[31-20] ^ c[31-21] ^ c[31-23] ^ c[31-25] ^ c[31-26] ^ c[31-28] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc512_crc[10] <= d[511-511] ^ d[511-510] ^ d[511-509] ^ d[511-507] ^ d[511-506] ^ d[511-504] ^ d[511-502] ^ d[511-501] ^ d[511-500] ^ d[511-499] ^ d[511-498] ^ d[511-494] ^ d[511-491] ^ d[511-488] ^ d[511-487] ^ d[511-484] ^ d[511-480] ^ d[511-479] ^ d[511-477] ^ d[511-471] ^ d[511-464] ^ d[511-463] ^ d[511-462] ^ d[511-460] ^ d[511-459] ^ d[511-457] ^ d[511-454] ^ d[511-449] ^ d[511-446] ^ d[511-445] ^ d[511-444] ^ d[511-442] ^ d[511-441] ^ d[511-438] ^ d[511-437] ^ d[511-436] ^ d[511-434] ^ d[511-432] ^ d[511-429] ^ d[511-428] ^ d[511-426] ^ d[511-425] ^ d[511-421] ^ d[511-420] ^ d[511-419] ^ d[511-418] ^ d[511-417] ^ d[511-416] ^ d[511-415] ^ d[511-413] ^ d[511-412] ^ d[511-411] ^ d[511-410] ^ d[511-409] ^ d[511-401] ^ d[511-400] ^ d[511-398] ^ d[511-397] ^ d[511-394] ^ d[511-392] ^ d[511-391] ^ d[511-389] ^ d[511-388] ^ d[511-387] ^ d[511-386] ^ d[511-384] ^ d[511-383] ^ d[511-376] ^ d[511-374] ^ d[511-372] ^ d[511-369] ^ d[511-368] ^ d[511-366] ^ d[511-362] ^ d[511-360] ^ d[511-358] ^ d[511-354] ^ d[511-353] ^ d[511-352] ^ d[511-348] ^ d[511-347] ^ d[511-346] ^ d[511-345] ^ d[511-343] ^ d[511-342] ^ d[511-341] ^ d[511-340] ^ d[511-335] ^ d[511-334] ^ d[511-332] ^ d[511-329] ^ d[511-326] ^ d[511-325] ^ d[511-324] ^ d[511-321] ^ d[511-312] ^ d[511-310] ^ d[511-308] ^ d[511-307] ^ d[511-306] ^ d[511-305] ^ d[511-304] ^ d[511-303] ^ d[511-302] ^ d[511-301] ^ d[511-297] ^ d[511-295] ^ d[511-293] ^ d[511-292] ^ d[511-291] ^ d[511-289] ^ d[511-287] ^ d[511-286] ^ d[511-281] ^ d[511-279] ^ d[511-275] ^ d[511-273] ^ d[511-269] ^ d[511-268] ^ d[511-265] ^ d[511-255] ^ d[511-254] ^ d[511-252] ^ d[511-251] ^ d[511-250] ^ d[511-248] ^ d[511-244] ^ d[511-243] ^ d[511-242] ^ d[511-238] ^ d[511-237] ^ d[511-236] ^ d[511-235] ^ d[511-233] ^ d[511-232] ^ d[511-228] ^ d[511-227] ^ d[511-226] ^ d[511-225] ^ d[511-224] ^ d[511-223] ^ d[511-221] ^ d[511-217] ^ d[511-216] ^ d[511-214] ^ d[511-212] ^ d[511-210] ^ d[511-207] ^ d[511-205] ^ d[511-204] ^ d[511-201] ^ d[511-198] ^ d[511-195] ^ d[511-194] ^ d[511-191] ^ d[511-190] ^ d[511-189] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-184] ^ d[511-179] ^ d[511-178] ^ d[511-175] ^ d[511-172] ^ d[511-165] ^ d[511-162] ^ d[511-161] ^ d[511-160] ^ d[511-158] ^ d[511-156] ^ d[511-150] ^ d[511-149] ^ d[511-148] ^ d[511-146] ^ d[511-145] ^ d[511-143] ^ d[511-141] ^ d[511-140] ^ d[511-139] ^ d[511-136] ^ d[511-133] ^ d[511-132] ^ d[511-129] ^ d[511-126] ^ d[511-125] ^ d[511-124] ^ d[511-123] ^ d[511-121] ^ d[511-120] ^ d[511-117] ^ d[511-116] ^ d[511-115] ^ d[511-114] ^ d[511-110] ^ d[511-109] ^ d[511-108] ^ d[511-107] ^ d[511-105] ^ d[511-104] ^ d[511-102] ^ d[511-99] ^ d[511-96] ^ d[511-95] ^ d[511-94] ^ d[511-92] ^ d[511-91] ^ d[511-89] ^ d[511-88] ^ d[511-87] ^ d[511-83] ^ d[511-82] ^ d[511-80] ^ d[511-73] ^ d[511-71] ^ d[511-62] ^ d[511-61] ^ d[511-56] ^ d[511-53] ^ d[511-52] ^ d[511-51] ^ d[511-49] ^ d[511-42] ^ d[511-40] ^ d[511-37] ^ d[511-35] ^ d[511-34] ^ d[511-31] ^ d[511-29] ^ d[511-27] ^ d[511-26] ^ d[511-24] ^ d[511-22] ^ d[511-18] ^ d[511-17] ^ d[511-13] ^ d[511-10] ^ d[511-9] ^ d[511-5] ^ c[31-0] ^ c[31-4] ^ c[31-7] ^ c[31-8] ^ c[31-11] ^ c[31-14] ^ c[31-18] ^ c[31-19] ^ c[31-20] ^ c[31-21] ^ c[31-22] ^ c[31-24] ^ c[31-26] ^ c[31-27] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc512_crc[9] <= d[511-506] ^ d[511-505] ^ d[511-503] ^ d[511-499] ^ d[511-494] ^ d[511-493] ^ d[511-491] ^ d[511-490] ^ d[511-486] ^ d[511-485] ^ d[511-483] ^ d[511-482] ^ d[511-479] ^ d[511-478] ^ d[511-477] ^ d[511-476] ^ d[511-470] ^ d[511-468] ^ d[511-463] ^ d[511-462] ^ d[511-460] ^ d[511-455] ^ d[511-452] ^ d[511-449] ^ d[511-448] ^ d[511-447] ^ d[511-446] ^ d[511-445] ^ d[511-444] ^ d[511-443] ^ d[511-442] ^ d[511-439] ^ d[511-438] ^ d[511-436] ^ d[511-435] ^ d[511-434] ^ d[511-430] ^ d[511-429] ^ d[511-427] ^ d[511-426] ^ d[511-424] ^ d[511-421] ^ d[511-420] ^ d[511-417] ^ d[511-413] ^ d[511-411] ^ d[511-410] ^ d[511-409] ^ d[511-408] ^ d[511-407] ^ d[511-405] ^ d[511-404] ^ d[511-402] ^ d[511-401] ^ d[511-400] ^ d[511-396] ^ d[511-395] ^ d[511-391] ^ d[511-389] ^ d[511-386] ^ d[511-385] ^ d[511-384] ^ d[511-381] ^ d[511-378] ^ d[511-377] ^ d[511-376] ^ d[511-375] ^ d[511-374] ^ d[511-373] ^ d[511-372] ^ d[511-370] ^ d[511-368] ^ d[511-367] ^ d[511-366] ^ d[511-362] ^ d[511-361] ^ d[511-358] ^ d[511-357] ^ d[511-355] ^ d[511-354] ^ d[511-346] ^ d[511-345] ^ d[511-343] ^ d[511-339] ^ d[511-338] ^ d[511-337] ^ d[511-336] ^ d[511-334] ^ d[511-330] ^ d[511-328] ^ d[511-326] ^ d[511-325] ^ d[511-321] ^ d[511-320] ^ d[511-319] ^ d[511-318] ^ d[511-317] ^ d[511-315] ^ d[511-313] ^ d[511-312] ^ d[511-311] ^ d[511-310] ^ d[511-308] ^ d[511-307] ^ d[511-306] ^ d[511-304] ^ d[511-300] ^ d[511-299] ^ d[511-297] ^ d[511-295] ^ d[511-293] ^ d[511-286] ^ d[511-283] ^ d[511-282] ^ d[511-280] ^ d[511-279] ^ d[511-277] ^ d[511-273] ^ d[511-270] ^ d[511-268] ^ d[511-266] ^ d[511-265] ^ d[511-264] ^ d[511-261] ^ d[511-259] ^ d[511-257] ^ d[511-256] ^ d[511-253] ^ d[511-251] ^ d[511-249] ^ d[511-248] ^ d[511-245] ^ d[511-244] ^ d[511-239] ^ d[511-238] ^ d[511-236] ^ d[511-233] ^ d[511-230] ^ d[511-229] ^ d[511-225] ^ d[511-222] ^ d[511-218] ^ d[511-217] ^ d[511-216] ^ d[511-215] ^ d[511-214] ^ d[511-213] ^ d[511-212] ^ d[511-211] ^ d[511-210] ^ d[511-209] ^ d[511-207] ^ d[511-206] ^ d[511-205] ^ d[511-203] ^ d[511-201] ^ d[511-198] ^ d[511-197] ^ d[511-196] ^ d[511-195] ^ d[511-194] ^ d[511-193] ^ d[511-189] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-183] ^ d[511-182] ^ d[511-180] ^ d[511-179] ^ d[511-176] ^ d[511-173] ^ d[511-172] ^ d[511-171] ^ d[511-170] ^ d[511-169] ^ d[511-167] ^ d[511-163] ^ d[511-159] ^ d[511-158] ^ d[511-157] ^ d[511-156] ^ d[511-155] ^ d[511-150] ^ d[511-147] ^ d[511-146] ^ d[511-143] ^ d[511-142] ^ d[511-141] ^ d[511-140] ^ d[511-136] ^ d[511-135] ^ d[511-133] ^ d[511-132] ^ d[511-130] ^ d[511-128] ^ d[511-124] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-119] ^ d[511-115] ^ d[511-114] ^ d[511-113] ^ d[511-109] ^ d[511-108] ^ d[511-105] ^ d[511-104] ^ d[511-101] ^ d[511-100] ^ d[511-99] ^ d[511-98] ^ d[511-94] ^ d[511-93] ^ d[511-92] ^ d[511-90] ^ d[511-89] ^ d[511-88] ^ d[511-87] ^ d[511-85] ^ d[511-82] ^ d[511-79] ^ d[511-74] ^ d[511-73] ^ d[511-68] ^ d[511-67] ^ d[511-66] ^ d[511-65] ^ d[511-62] ^ d[511-61] ^ d[511-60] ^ d[511-58] ^ d[511-57] ^ d[511-55] ^ d[511-52] ^ d[511-48] ^ d[511-47] ^ d[511-45] ^ d[511-44] ^ d[511-43] ^ d[511-41] ^ d[511-38] ^ d[511-37] ^ d[511-36] ^ d[511-35] ^ d[511-34] ^ d[511-31] ^ d[511-29] ^ d[511-27] ^ d[511-26] ^ d[511-24] ^ d[511-23] ^ d[511-19] ^ d[511-18] ^ d[511-16] ^ d[511-14] ^ d[511-12] ^ d[511-11] ^ d[511-9] ^ d[511-0] ^ c[31-2] ^ c[31-3] ^ c[31-5] ^ c[31-6] ^ c[31-10] ^ c[31-11] ^ c[31-13] ^ c[31-14] ^ c[31-19] ^ c[31-23] ^ c[31-25] ^ c[31-26];
                stage_crc512_crc[8] <= d[511-511] ^ d[511-510] ^ d[511-508] ^ d[511-504] ^ d[511-502] ^ d[511-501] ^ d[511-493] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-487] ^ d[511-484] ^ d[511-482] ^ d[511-481] ^ d[511-478] ^ d[511-476] ^ d[511-472] ^ d[511-471] ^ d[511-470] ^ d[511-469] ^ d[511-468] ^ d[511-465] ^ d[511-463] ^ d[511-462] ^ d[511-458] ^ d[511-456] ^ d[511-453] ^ d[511-452] ^ d[511-447] ^ d[511-446] ^ d[511-445] ^ d[511-443] ^ d[511-440] ^ d[511-439] ^ d[511-435] ^ d[511-434] ^ d[511-433] ^ d[511-431] ^ d[511-430] ^ d[511-428] ^ d[511-427] ^ d[511-425] ^ d[511-424] ^ d[511-421] ^ d[511-419] ^ d[511-416] ^ d[511-411] ^ d[511-410] ^ d[511-407] ^ d[511-406] ^ d[511-404] ^ d[511-403] ^ d[511-402] ^ d[511-401] ^ d[511-400] ^ d[511-399] ^ d[511-398] ^ d[511-397] ^ d[511-393] ^ d[511-391] ^ d[511-388] ^ d[511-385] ^ d[511-382] ^ d[511-381] ^ d[511-379] ^ d[511-377] ^ d[511-375] ^ d[511-373] ^ d[511-372] ^ d[511-371] ^ d[511-367] ^ d[511-366] ^ d[511-357] ^ d[511-356] ^ d[511-355] ^ d[511-353] ^ d[511-349] ^ d[511-348] ^ d[511-346] ^ d[511-345] ^ d[511-342] ^ d[511-341] ^ d[511-340] ^ d[511-334] ^ d[511-333] ^ d[511-331] ^ d[511-329] ^ d[511-328] ^ d[511-326] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-313] ^ d[511-311] ^ d[511-310] ^ d[511-308] ^ d[511-307] ^ d[511-303] ^ d[511-302] ^ d[511-301] ^ d[511-299] ^ d[511-297] ^ d[511-295] ^ d[511-292] ^ d[511-290] ^ d[511-288] ^ d[511-286] ^ d[511-284] ^ d[511-281] ^ d[511-280] ^ d[511-279] ^ d[511-278] ^ d[511-277] ^ d[511-276] ^ d[511-273] ^ d[511-271] ^ d[511-268] ^ d[511-267] ^ d[511-266] ^ d[511-264] ^ d[511-262] ^ d[511-261] ^ d[511-260] ^ d[511-259] ^ d[511-258] ^ d[511-255] ^ d[511-254] ^ d[511-250] ^ d[511-249] ^ d[511-248] ^ d[511-246] ^ d[511-245] ^ d[511-243] ^ d[511-240] ^ d[511-239] ^ d[511-231] ^ d[511-228] ^ d[511-227] ^ d[511-224] ^ d[511-223] ^ d[511-219] ^ d[511-218] ^ d[511-217] ^ d[511-215] ^ d[511-213] ^ d[511-211] ^ d[511-209] ^ d[511-206] ^ d[511-204] ^ d[511-203] ^ d[511-201] ^ d[511-196] ^ d[511-195] ^ d[511-193] ^ d[511-192] ^ d[511-191] ^ d[511-187] ^ d[511-184] ^ d[511-182] ^ d[511-181] ^ d[511-180] ^ d[511-177] ^ d[511-174] ^ d[511-173] ^ d[511-169] ^ d[511-168] ^ d[511-167] ^ d[511-166] ^ d[511-164] ^ d[511-162] ^ d[511-161] ^ d[511-160] ^ d[511-159] ^ d[511-157] ^ d[511-155] ^ d[511-149] ^ d[511-148] ^ d[511-147] ^ d[511-142] ^ d[511-141] ^ d[511-135] ^ d[511-133] ^ d[511-132] ^ d[511-131] ^ d[511-129] ^ d[511-128] ^ d[511-127] ^ d[511-126] ^ d[511-124] ^ d[511-122] ^ d[511-120] ^ d[511-119] ^ d[511-118] ^ d[511-117] ^ d[511-115] ^ d[511-113] ^ d[511-111] ^ d[511-109] ^ d[511-105] ^ d[511-104] ^ d[511-103] ^ d[511-102] ^ d[511-100] ^ d[511-98] ^ d[511-97] ^ d[511-96] ^ d[511-93] ^ d[511-91] ^ d[511-90] ^ d[511-89] ^ d[511-88] ^ d[511-87] ^ d[511-86] ^ d[511-85] ^ d[511-84] ^ d[511-82] ^ d[511-81] ^ d[511-80] ^ d[511-79] ^ d[511-75] ^ d[511-74] ^ d[511-73] ^ d[511-72] ^ d[511-69] ^ d[511-65] ^ d[511-62] ^ d[511-60] ^ d[511-59] ^ d[511-56] ^ d[511-55] ^ d[511-54] ^ d[511-50] ^ d[511-49] ^ d[511-47] ^ d[511-46] ^ d[511-42] ^ d[511-39] ^ d[511-38] ^ d[511-36] ^ d[511-35] ^ d[511-34] ^ d[511-31] ^ d[511-29] ^ d[511-27] ^ d[511-26] ^ d[511-20] ^ d[511-19] ^ d[511-17] ^ d[511-16] ^ d[511-15] ^ d[511-13] ^ d[511-9] ^ d[511-6] ^ d[511-1] ^ d[511-0] ^ c[31-1] ^ c[31-2] ^ c[31-4] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-13] ^ c[31-21] ^ c[31-22] ^ c[31-24] ^ c[31-28] ^ c[31-30] ^ c[31-31];
                stage_crc512_crc[7] <= d[511-511] ^ d[511-509] ^ d[511-505] ^ d[511-503] ^ d[511-502] ^ d[511-494] ^ d[511-491] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-485] ^ d[511-483] ^ d[511-482] ^ d[511-479] ^ d[511-477] ^ d[511-473] ^ d[511-472] ^ d[511-471] ^ d[511-470] ^ d[511-469] ^ d[511-466] ^ d[511-464] ^ d[511-463] ^ d[511-459] ^ d[511-457] ^ d[511-454] ^ d[511-453] ^ d[511-448] ^ d[511-447] ^ d[511-446] ^ d[511-444] ^ d[511-441] ^ d[511-440] ^ d[511-436] ^ d[511-435] ^ d[511-434] ^ d[511-432] ^ d[511-431] ^ d[511-429] ^ d[511-428] ^ d[511-426] ^ d[511-425] ^ d[511-422] ^ d[511-420] ^ d[511-417] ^ d[511-412] ^ d[511-411] ^ d[511-408] ^ d[511-407] ^ d[511-405] ^ d[511-404] ^ d[511-403] ^ d[511-402] ^ d[511-401] ^ d[511-400] ^ d[511-399] ^ d[511-398] ^ d[511-394] ^ d[511-392] ^ d[511-389] ^ d[511-386] ^ d[511-383] ^ d[511-382] ^ d[511-380] ^ d[511-378] ^ d[511-376] ^ d[511-374] ^ d[511-373] ^ d[511-372] ^ d[511-368] ^ d[511-367] ^ d[511-358] ^ d[511-357] ^ d[511-356] ^ d[511-354] ^ d[511-350] ^ d[511-349] ^ d[511-347] ^ d[511-346] ^ d[511-343] ^ d[511-342] ^ d[511-341] ^ d[511-335] ^ d[511-334] ^ d[511-332] ^ d[511-330] ^ d[511-329] ^ d[511-327] ^ d[511-318] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-312] ^ d[511-311] ^ d[511-309] ^ d[511-308] ^ d[511-304] ^ d[511-303] ^ d[511-302] ^ d[511-300] ^ d[511-298] ^ d[511-296] ^ d[511-293] ^ d[511-291] ^ d[511-289] ^ d[511-287] ^ d[511-285] ^ d[511-282] ^ d[511-281] ^ d[511-280] ^ d[511-279] ^ d[511-278] ^ d[511-277] ^ d[511-274] ^ d[511-272] ^ d[511-269] ^ d[511-268] ^ d[511-267] ^ d[511-265] ^ d[511-263] ^ d[511-262] ^ d[511-261] ^ d[511-260] ^ d[511-259] ^ d[511-256] ^ d[511-255] ^ d[511-251] ^ d[511-250] ^ d[511-249] ^ d[511-247] ^ d[511-246] ^ d[511-244] ^ d[511-241] ^ d[511-240] ^ d[511-232] ^ d[511-229] ^ d[511-228] ^ d[511-225] ^ d[511-224] ^ d[511-220] ^ d[511-219] ^ d[511-218] ^ d[511-216] ^ d[511-214] ^ d[511-212] ^ d[511-210] ^ d[511-207] ^ d[511-205] ^ d[511-204] ^ d[511-202] ^ d[511-197] ^ d[511-196] ^ d[511-194] ^ d[511-193] ^ d[511-192] ^ d[511-188] ^ d[511-185] ^ d[511-183] ^ d[511-182] ^ d[511-181] ^ d[511-178] ^ d[511-175] ^ d[511-174] ^ d[511-170] ^ d[511-169] ^ d[511-168] ^ d[511-167] ^ d[511-165] ^ d[511-163] ^ d[511-162] ^ d[511-161] ^ d[511-160] ^ d[511-158] ^ d[511-156] ^ d[511-150] ^ d[511-149] ^ d[511-148] ^ d[511-143] ^ d[511-142] ^ d[511-136] ^ d[511-134] ^ d[511-133] ^ d[511-132] ^ d[511-130] ^ d[511-129] ^ d[511-128] ^ d[511-127] ^ d[511-125] ^ d[511-123] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-118] ^ d[511-116] ^ d[511-114] ^ d[511-112] ^ d[511-110] ^ d[511-106] ^ d[511-105] ^ d[511-104] ^ d[511-103] ^ d[511-101] ^ d[511-99] ^ d[511-98] ^ d[511-97] ^ d[511-94] ^ d[511-92] ^ d[511-91] ^ d[511-90] ^ d[511-89] ^ d[511-88] ^ d[511-87] ^ d[511-86] ^ d[511-85] ^ d[511-83] ^ d[511-82] ^ d[511-81] ^ d[511-80] ^ d[511-76] ^ d[511-75] ^ d[511-74] ^ d[511-73] ^ d[511-70] ^ d[511-66] ^ d[511-63] ^ d[511-61] ^ d[511-60] ^ d[511-57] ^ d[511-56] ^ d[511-55] ^ d[511-51] ^ d[511-50] ^ d[511-48] ^ d[511-47] ^ d[511-43] ^ d[511-40] ^ d[511-39] ^ d[511-37] ^ d[511-36] ^ d[511-35] ^ d[511-32] ^ d[511-30] ^ d[511-28] ^ d[511-27] ^ d[511-21] ^ d[511-20] ^ d[511-18] ^ d[511-17] ^ d[511-16] ^ d[511-14] ^ d[511-10] ^ d[511-7] ^ d[511-2] ^ d[511-1] ^ c[31-2] ^ c[31-3] ^ c[31-5] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-14] ^ c[31-22] ^ c[31-23] ^ c[31-25] ^ c[31-29] ^ c[31-31];
                stage_crc512_crc[6] <= d[511-510] ^ d[511-506] ^ d[511-504] ^ d[511-503] ^ d[511-495] ^ d[511-492] ^ d[511-491] ^ d[511-490] ^ d[511-489] ^ d[511-486] ^ d[511-484] ^ d[511-483] ^ d[511-480] ^ d[511-478] ^ d[511-474] ^ d[511-473] ^ d[511-472] ^ d[511-471] ^ d[511-470] ^ d[511-467] ^ d[511-465] ^ d[511-464] ^ d[511-460] ^ d[511-458] ^ d[511-455] ^ d[511-454] ^ d[511-449] ^ d[511-448] ^ d[511-447] ^ d[511-445] ^ d[511-442] ^ d[511-441] ^ d[511-437] ^ d[511-436] ^ d[511-435] ^ d[511-433] ^ d[511-432] ^ d[511-430] ^ d[511-429] ^ d[511-427] ^ d[511-426] ^ d[511-423] ^ d[511-421] ^ d[511-418] ^ d[511-413] ^ d[511-412] ^ d[511-409] ^ d[511-408] ^ d[511-406] ^ d[511-405] ^ d[511-404] ^ d[511-403] ^ d[511-402] ^ d[511-401] ^ d[511-400] ^ d[511-399] ^ d[511-395] ^ d[511-393] ^ d[511-390] ^ d[511-387] ^ d[511-384] ^ d[511-383] ^ d[511-381] ^ d[511-379] ^ d[511-377] ^ d[511-375] ^ d[511-374] ^ d[511-373] ^ d[511-369] ^ d[511-368] ^ d[511-359] ^ d[511-358] ^ d[511-357] ^ d[511-355] ^ d[511-351] ^ d[511-350] ^ d[511-348] ^ d[511-347] ^ d[511-344] ^ d[511-343] ^ d[511-342] ^ d[511-336] ^ d[511-335] ^ d[511-333] ^ d[511-331] ^ d[511-330] ^ d[511-328] ^ d[511-319] ^ d[511-318] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-313] ^ d[511-312] ^ d[511-310] ^ d[511-309] ^ d[511-305] ^ d[511-304] ^ d[511-303] ^ d[511-301] ^ d[511-299] ^ d[511-297] ^ d[511-294] ^ d[511-292] ^ d[511-290] ^ d[511-288] ^ d[511-286] ^ d[511-283] ^ d[511-282] ^ d[511-281] ^ d[511-280] ^ d[511-279] ^ d[511-278] ^ d[511-275] ^ d[511-273] ^ d[511-270] ^ d[511-269] ^ d[511-268] ^ d[511-266] ^ d[511-264] ^ d[511-263] ^ d[511-262] ^ d[511-261] ^ d[511-260] ^ d[511-257] ^ d[511-256] ^ d[511-252] ^ d[511-251] ^ d[511-250] ^ d[511-248] ^ d[511-247] ^ d[511-245] ^ d[511-242] ^ d[511-241] ^ d[511-233] ^ d[511-230] ^ d[511-229] ^ d[511-226] ^ d[511-225] ^ d[511-221] ^ d[511-220] ^ d[511-219] ^ d[511-217] ^ d[511-215] ^ d[511-213] ^ d[511-211] ^ d[511-208] ^ d[511-206] ^ d[511-205] ^ d[511-203] ^ d[511-198] ^ d[511-197] ^ d[511-195] ^ d[511-194] ^ d[511-193] ^ d[511-189] ^ d[511-186] ^ d[511-184] ^ d[511-183] ^ d[511-182] ^ d[511-179] ^ d[511-176] ^ d[511-175] ^ d[511-171] ^ d[511-170] ^ d[511-169] ^ d[511-168] ^ d[511-166] ^ d[511-164] ^ d[511-163] ^ d[511-162] ^ d[511-161] ^ d[511-159] ^ d[511-157] ^ d[511-151] ^ d[511-150] ^ d[511-149] ^ d[511-144] ^ d[511-143] ^ d[511-137] ^ d[511-135] ^ d[511-134] ^ d[511-133] ^ d[511-131] ^ d[511-130] ^ d[511-129] ^ d[511-128] ^ d[511-126] ^ d[511-124] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-117] ^ d[511-115] ^ d[511-113] ^ d[511-111] ^ d[511-107] ^ d[511-106] ^ d[511-105] ^ d[511-104] ^ d[511-102] ^ d[511-100] ^ d[511-99] ^ d[511-98] ^ d[511-95] ^ d[511-93] ^ d[511-92] ^ d[511-91] ^ d[511-90] ^ d[511-89] ^ d[511-88] ^ d[511-87] ^ d[511-86] ^ d[511-84] ^ d[511-83] ^ d[511-82] ^ d[511-81] ^ d[511-77] ^ d[511-76] ^ d[511-75] ^ d[511-74] ^ d[511-71] ^ d[511-67] ^ d[511-64] ^ d[511-62] ^ d[511-61] ^ d[511-58] ^ d[511-57] ^ d[511-56] ^ d[511-52] ^ d[511-51] ^ d[511-49] ^ d[511-48] ^ d[511-44] ^ d[511-41] ^ d[511-40] ^ d[511-38] ^ d[511-37] ^ d[511-36] ^ d[511-33] ^ d[511-31] ^ d[511-29] ^ d[511-28] ^ d[511-22] ^ d[511-21] ^ d[511-19] ^ d[511-18] ^ d[511-17] ^ d[511-15] ^ d[511-11] ^ d[511-8] ^ d[511-3] ^ d[511-2] ^ c[31-0] ^ c[31-3] ^ c[31-4] ^ c[31-6] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-15] ^ c[31-23] ^ c[31-24] ^ c[31-26] ^ c[31-30];
                stage_crc512_crc[5] <= d[511-510] ^ d[511-508] ^ d[511-506] ^ d[511-505] ^ d[511-504] ^ d[511-502] ^ d[511-501] ^ d[511-500] ^ d[511-496] ^ d[511-495] ^ d[511-494] ^ d[511-489] ^ d[511-488] ^ d[511-487] ^ d[511-486] ^ d[511-485] ^ d[511-484] ^ d[511-483] ^ d[511-482] ^ d[511-480] ^ d[511-477] ^ d[511-476] ^ d[511-475] ^ d[511-474] ^ d[511-473] ^ d[511-471] ^ d[511-470] ^ d[511-466] ^ d[511-464] ^ d[511-462] ^ d[511-459] ^ d[511-458] ^ d[511-456] ^ d[511-455] ^ d[511-452] ^ d[511-446] ^ d[511-444] ^ d[511-443] ^ d[511-442] ^ d[511-438] ^ d[511-431] ^ d[511-430] ^ d[511-428] ^ d[511-427] ^ d[511-418] ^ d[511-416] ^ d[511-413] ^ d[511-412] ^ d[511-410] ^ d[511-408] ^ d[511-406] ^ d[511-403] ^ d[511-402] ^ d[511-401] ^ d[511-399] ^ d[511-398] ^ d[511-394] ^ d[511-393] ^ d[511-392] ^ d[511-390] ^ d[511-387] ^ d[511-386] ^ d[511-385] ^ d[511-384] ^ d[511-382] ^ d[511-381] ^ d[511-380] ^ d[511-375] ^ d[511-372] ^ d[511-370] ^ d[511-368] ^ d[511-366] ^ d[511-363] ^ d[511-362] ^ d[511-360] ^ d[511-357] ^ d[511-356] ^ d[511-353] ^ d[511-352] ^ d[511-351] ^ d[511-347] ^ d[511-343] ^ d[511-342] ^ d[511-341] ^ d[511-339] ^ d[511-338] ^ d[511-336] ^ d[511-335] ^ d[511-333] ^ d[511-332] ^ d[511-331] ^ d[511-329] ^ d[511-328] ^ d[511-327] ^ d[511-322] ^ d[511-321] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-313] ^ d[511-312] ^ d[511-311] ^ d[511-309] ^ d[511-306] ^ d[511-304] ^ d[511-303] ^ d[511-299] ^ d[511-297] ^ d[511-296] ^ d[511-294] ^ d[511-293] ^ d[511-292] ^ d[511-291] ^ d[511-290] ^ d[511-289] ^ d[511-288] ^ d[511-286] ^ d[511-284] ^ d[511-282] ^ d[511-281] ^ d[511-280] ^ d[511-277] ^ d[511-273] ^ d[511-271] ^ d[511-270] ^ d[511-268] ^ d[511-267] ^ d[511-263] ^ d[511-262] ^ d[511-259] ^ d[511-258] ^ d[511-255] ^ d[511-253] ^ d[511-251] ^ d[511-249] ^ d[511-246] ^ d[511-242] ^ d[511-237] ^ d[511-231] ^ d[511-228] ^ d[511-224] ^ d[511-222] ^ d[511-221] ^ d[511-220] ^ d[511-218] ^ d[511-210] ^ d[511-208] ^ d[511-206] ^ d[511-204] ^ d[511-203] ^ d[511-202] ^ d[511-201] ^ d[511-197] ^ d[511-196] ^ d[511-195] ^ d[511-193] ^ d[511-192] ^ d[511-191] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-184] ^ d[511-182] ^ d[511-180] ^ d[511-177] ^ d[511-176] ^ d[511-166] ^ d[511-165] ^ d[511-164] ^ d[511-163] ^ d[511-161] ^ d[511-160] ^ d[511-156] ^ d[511-155] ^ d[511-152] ^ d[511-150] ^ d[511-149] ^ d[511-145] ^ d[511-143] ^ d[511-138] ^ d[511-137] ^ d[511-131] ^ d[511-130] ^ d[511-129] ^ d[511-128] ^ d[511-126] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-119] ^ d[511-117] ^ d[511-113] ^ d[511-112] ^ d[511-111] ^ d[511-110] ^ d[511-108] ^ d[511-107] ^ d[511-105] ^ d[511-104] ^ d[511-100] ^ d[511-98] ^ d[511-97] ^ d[511-95] ^ d[511-93] ^ d[511-92] ^ d[511-91] ^ d[511-90] ^ d[511-89] ^ d[511-88] ^ d[511-81] ^ d[511-79] ^ d[511-78] ^ d[511-77] ^ d[511-76] ^ d[511-75] ^ d[511-73] ^ d[511-67] ^ d[511-66] ^ d[511-62] ^ d[511-61] ^ d[511-60] ^ d[511-59] ^ d[511-57] ^ d[511-55] ^ d[511-54] ^ d[511-52] ^ d[511-49] ^ d[511-48] ^ d[511-47] ^ d[511-44] ^ d[511-42] ^ d[511-41] ^ d[511-39] ^ d[511-38] ^ d[511-31] ^ d[511-28] ^ d[511-26] ^ d[511-25] ^ d[511-24] ^ d[511-23] ^ d[511-22] ^ d[511-20] ^ d[511-19] ^ d[511-18] ^ d[511-10] ^ d[511-6] ^ d[511-4] ^ d[511-3] ^ d[511-0] ^ c[31-0] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-20] ^ c[31-21] ^ c[31-22] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-28] ^ c[31-30];
                stage_crc512_crc[4] <= d[511-511] ^ d[511-509] ^ d[511-507] ^ d[511-506] ^ d[511-505] ^ d[511-503] ^ d[511-502] ^ d[511-501] ^ d[511-497] ^ d[511-496] ^ d[511-495] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-487] ^ d[511-486] ^ d[511-485] ^ d[511-484] ^ d[511-483] ^ d[511-481] ^ d[511-478] ^ d[511-477] ^ d[511-476] ^ d[511-475] ^ d[511-474] ^ d[511-472] ^ d[511-471] ^ d[511-467] ^ d[511-465] ^ d[511-463] ^ d[511-460] ^ d[511-459] ^ d[511-457] ^ d[511-456] ^ d[511-453] ^ d[511-447] ^ d[511-445] ^ d[511-444] ^ d[511-443] ^ d[511-439] ^ d[511-432] ^ d[511-431] ^ d[511-429] ^ d[511-428] ^ d[511-419] ^ d[511-417] ^ d[511-414] ^ d[511-413] ^ d[511-411] ^ d[511-409] ^ d[511-407] ^ d[511-404] ^ d[511-403] ^ d[511-402] ^ d[511-400] ^ d[511-399] ^ d[511-395] ^ d[511-394] ^ d[511-393] ^ d[511-391] ^ d[511-388] ^ d[511-387] ^ d[511-386] ^ d[511-385] ^ d[511-383] ^ d[511-382] ^ d[511-381] ^ d[511-376] ^ d[511-373] ^ d[511-371] ^ d[511-369] ^ d[511-367] ^ d[511-364] ^ d[511-363] ^ d[511-361] ^ d[511-358] ^ d[511-357] ^ d[511-354] ^ d[511-353] ^ d[511-352] ^ d[511-348] ^ d[511-344] ^ d[511-343] ^ d[511-342] ^ d[511-340] ^ d[511-339] ^ d[511-337] ^ d[511-336] ^ d[511-334] ^ d[511-333] ^ d[511-332] ^ d[511-330] ^ d[511-329] ^ d[511-328] ^ d[511-323] ^ d[511-322] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-313] ^ d[511-312] ^ d[511-310] ^ d[511-307] ^ d[511-305] ^ d[511-304] ^ d[511-300] ^ d[511-298] ^ d[511-297] ^ d[511-295] ^ d[511-294] ^ d[511-293] ^ d[511-292] ^ d[511-291] ^ d[511-290] ^ d[511-289] ^ d[511-287] ^ d[511-285] ^ d[511-283] ^ d[511-282] ^ d[511-281] ^ d[511-278] ^ d[511-274] ^ d[511-272] ^ d[511-271] ^ d[511-269] ^ d[511-268] ^ d[511-264] ^ d[511-263] ^ d[511-260] ^ d[511-259] ^ d[511-256] ^ d[511-254] ^ d[511-252] ^ d[511-250] ^ d[511-247] ^ d[511-243] ^ d[511-238] ^ d[511-232] ^ d[511-229] ^ d[511-225] ^ d[511-223] ^ d[511-222] ^ d[511-221] ^ d[511-219] ^ d[511-211] ^ d[511-209] ^ d[511-207] ^ d[511-205] ^ d[511-204] ^ d[511-203] ^ d[511-202] ^ d[511-198] ^ d[511-197] ^ d[511-196] ^ d[511-194] ^ d[511-193] ^ d[511-192] ^ d[511-189] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-185] ^ d[511-183] ^ d[511-181] ^ d[511-178] ^ d[511-177] ^ d[511-167] ^ d[511-166] ^ d[511-165] ^ d[511-164] ^ d[511-162] ^ d[511-161] ^ d[511-157] ^ d[511-156] ^ d[511-153] ^ d[511-151] ^ d[511-150] ^ d[511-146] ^ d[511-144] ^ d[511-139] ^ d[511-138] ^ d[511-132] ^ d[511-131] ^ d[511-130] ^ d[511-129] ^ d[511-127] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-120] ^ d[511-118] ^ d[511-114] ^ d[511-113] ^ d[511-112] ^ d[511-111] ^ d[511-109] ^ d[511-108] ^ d[511-106] ^ d[511-105] ^ d[511-101] ^ d[511-99] ^ d[511-98] ^ d[511-96] ^ d[511-94] ^ d[511-93] ^ d[511-92] ^ d[511-91] ^ d[511-90] ^ d[511-89] ^ d[511-82] ^ d[511-80] ^ d[511-79] ^ d[511-78] ^ d[511-77] ^ d[511-76] ^ d[511-74] ^ d[511-68] ^ d[511-67] ^ d[511-63] ^ d[511-62] ^ d[511-61] ^ d[511-60] ^ d[511-58] ^ d[511-56] ^ d[511-55] ^ d[511-53] ^ d[511-50] ^ d[511-49] ^ d[511-48] ^ d[511-45] ^ d[511-43] ^ d[511-42] ^ d[511-40] ^ d[511-39] ^ d[511-32] ^ d[511-29] ^ d[511-27] ^ d[511-26] ^ d[511-25] ^ d[511-24] ^ d[511-23] ^ d[511-21] ^ d[511-20] ^ d[511-19] ^ d[511-11] ^ d[511-7] ^ d[511-5] ^ d[511-4] ^ d[511-1] ^ c[31-1] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-21] ^ c[31-22] ^ c[31-23] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-29] ^ c[31-31];
                stage_crc512_crc[3] <= d[511-510] ^ d[511-508] ^ d[511-507] ^ d[511-506] ^ d[511-504] ^ d[511-503] ^ d[511-502] ^ d[511-498] ^ d[511-497] ^ d[511-496] ^ d[511-491] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-487] ^ d[511-486] ^ d[511-485] ^ d[511-484] ^ d[511-482] ^ d[511-479] ^ d[511-478] ^ d[511-477] ^ d[511-476] ^ d[511-475] ^ d[511-473] ^ d[511-472] ^ d[511-468] ^ d[511-466] ^ d[511-464] ^ d[511-461] ^ d[511-460] ^ d[511-458] ^ d[511-457] ^ d[511-454] ^ d[511-448] ^ d[511-446] ^ d[511-445] ^ d[511-444] ^ d[511-440] ^ d[511-433] ^ d[511-432] ^ d[511-430] ^ d[511-429] ^ d[511-420] ^ d[511-418] ^ d[511-415] ^ d[511-414] ^ d[511-412] ^ d[511-410] ^ d[511-408] ^ d[511-405] ^ d[511-404] ^ d[511-403] ^ d[511-401] ^ d[511-400] ^ d[511-396] ^ d[511-395] ^ d[511-394] ^ d[511-392] ^ d[511-389] ^ d[511-388] ^ d[511-387] ^ d[511-386] ^ d[511-384] ^ d[511-383] ^ d[511-382] ^ d[511-377] ^ d[511-374] ^ d[511-372] ^ d[511-370] ^ d[511-368] ^ d[511-365] ^ d[511-364] ^ d[511-362] ^ d[511-359] ^ d[511-358] ^ d[511-355] ^ d[511-354] ^ d[511-353] ^ d[511-349] ^ d[511-345] ^ d[511-344] ^ d[511-343] ^ d[511-341] ^ d[511-340] ^ d[511-338] ^ d[511-337] ^ d[511-335] ^ d[511-334] ^ d[511-333] ^ d[511-331] ^ d[511-330] ^ d[511-329] ^ d[511-324] ^ d[511-323] ^ d[511-318] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-313] ^ d[511-311] ^ d[511-308] ^ d[511-306] ^ d[511-305] ^ d[511-301] ^ d[511-299] ^ d[511-298] ^ d[511-296] ^ d[511-295] ^ d[511-294] ^ d[511-293] ^ d[511-292] ^ d[511-291] ^ d[511-290] ^ d[511-288] ^ d[511-286] ^ d[511-284] ^ d[511-283] ^ d[511-282] ^ d[511-279] ^ d[511-275] ^ d[511-273] ^ d[511-272] ^ d[511-270] ^ d[511-269] ^ d[511-265] ^ d[511-264] ^ d[511-261] ^ d[511-260] ^ d[511-257] ^ d[511-255] ^ d[511-253] ^ d[511-251] ^ d[511-248] ^ d[511-244] ^ d[511-239] ^ d[511-233] ^ d[511-230] ^ d[511-226] ^ d[511-224] ^ d[511-223] ^ d[511-222] ^ d[511-220] ^ d[511-212] ^ d[511-210] ^ d[511-208] ^ d[511-206] ^ d[511-205] ^ d[511-204] ^ d[511-203] ^ d[511-199] ^ d[511-198] ^ d[511-197] ^ d[511-195] ^ d[511-194] ^ d[511-193] ^ d[511-190] ^ d[511-189] ^ d[511-188] ^ d[511-187] ^ d[511-186] ^ d[511-184] ^ d[511-182] ^ d[511-179] ^ d[511-178] ^ d[511-168] ^ d[511-167] ^ d[511-166] ^ d[511-165] ^ d[511-163] ^ d[511-162] ^ d[511-158] ^ d[511-157] ^ d[511-154] ^ d[511-152] ^ d[511-151] ^ d[511-147] ^ d[511-145] ^ d[511-140] ^ d[511-139] ^ d[511-133] ^ d[511-132] ^ d[511-131] ^ d[511-130] ^ d[511-128] ^ d[511-124] ^ d[511-123] ^ d[511-122] ^ d[511-121] ^ d[511-119] ^ d[511-115] ^ d[511-114] ^ d[511-113] ^ d[511-112] ^ d[511-110] ^ d[511-109] ^ d[511-107] ^ d[511-106] ^ d[511-102] ^ d[511-100] ^ d[511-99] ^ d[511-97] ^ d[511-95] ^ d[511-94] ^ d[511-93] ^ d[511-92] ^ d[511-91] ^ d[511-90] ^ d[511-83] ^ d[511-81] ^ d[511-80] ^ d[511-79] ^ d[511-78] ^ d[511-77] ^ d[511-75] ^ d[511-69] ^ d[511-68] ^ d[511-64] ^ d[511-63] ^ d[511-62] ^ d[511-61] ^ d[511-59] ^ d[511-57] ^ d[511-56] ^ d[511-54] ^ d[511-51] ^ d[511-50] ^ d[511-49] ^ d[511-46] ^ d[511-44] ^ d[511-43] ^ d[511-41] ^ d[511-40] ^ d[511-33] ^ d[511-30] ^ d[511-28] ^ d[511-27] ^ d[511-26] ^ d[511-25] ^ d[511-24] ^ d[511-22] ^ d[511-21] ^ d[511-20] ^ d[511-12] ^ d[511-8] ^ d[511-6] ^ d[511-5] ^ d[511-2] ^ c[31-2] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-22] ^ c[31-23] ^ c[31-24] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-30];
                stage_crc512_crc[2] <= d[511-511] ^ d[511-509] ^ d[511-508] ^ d[511-507] ^ d[511-505] ^ d[511-504] ^ d[511-503] ^ d[511-499] ^ d[511-498] ^ d[511-497] ^ d[511-492] ^ d[511-491] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-487] ^ d[511-486] ^ d[511-485] ^ d[511-483] ^ d[511-480] ^ d[511-479] ^ d[511-478] ^ d[511-477] ^ d[511-476] ^ d[511-474] ^ d[511-473] ^ d[511-469] ^ d[511-467] ^ d[511-465] ^ d[511-462] ^ d[511-461] ^ d[511-459] ^ d[511-458] ^ d[511-455] ^ d[511-449] ^ d[511-447] ^ d[511-446] ^ d[511-445] ^ d[511-441] ^ d[511-434] ^ d[511-433] ^ d[511-431] ^ d[511-430] ^ d[511-421] ^ d[511-419] ^ d[511-416] ^ d[511-415] ^ d[511-413] ^ d[511-411] ^ d[511-409] ^ d[511-406] ^ d[511-405] ^ d[511-404] ^ d[511-402] ^ d[511-401] ^ d[511-397] ^ d[511-396] ^ d[511-395] ^ d[511-393] ^ d[511-390] ^ d[511-389] ^ d[511-388] ^ d[511-387] ^ d[511-385] ^ d[511-384] ^ d[511-383] ^ d[511-378] ^ d[511-375] ^ d[511-373] ^ d[511-371] ^ d[511-369] ^ d[511-366] ^ d[511-365] ^ d[511-363] ^ d[511-360] ^ d[511-359] ^ d[511-356] ^ d[511-355] ^ d[511-354] ^ d[511-350] ^ d[511-346] ^ d[511-345] ^ d[511-344] ^ d[511-342] ^ d[511-341] ^ d[511-339] ^ d[511-338] ^ d[511-336] ^ d[511-335] ^ d[511-334] ^ d[511-332] ^ d[511-331] ^ d[511-330] ^ d[511-325] ^ d[511-324] ^ d[511-319] ^ d[511-318] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-314] ^ d[511-312] ^ d[511-309] ^ d[511-307] ^ d[511-306] ^ d[511-302] ^ d[511-300] ^ d[511-299] ^ d[511-297] ^ d[511-296] ^ d[511-295] ^ d[511-294] ^ d[511-293] ^ d[511-292] ^ d[511-291] ^ d[511-289] ^ d[511-287] ^ d[511-285] ^ d[511-284] ^ d[511-283] ^ d[511-280] ^ d[511-276] ^ d[511-274] ^ d[511-273] ^ d[511-271] ^ d[511-270] ^ d[511-266] ^ d[511-265] ^ d[511-262] ^ d[511-261] ^ d[511-258] ^ d[511-256] ^ d[511-254] ^ d[511-252] ^ d[511-249] ^ d[511-245] ^ d[511-240] ^ d[511-234] ^ d[511-231] ^ d[511-227] ^ d[511-225] ^ d[511-224] ^ d[511-223] ^ d[511-221] ^ d[511-213] ^ d[511-211] ^ d[511-209] ^ d[511-207] ^ d[511-206] ^ d[511-205] ^ d[511-204] ^ d[511-200] ^ d[511-199] ^ d[511-198] ^ d[511-196] ^ d[511-195] ^ d[511-194] ^ d[511-191] ^ d[511-190] ^ d[511-189] ^ d[511-188] ^ d[511-187] ^ d[511-185] ^ d[511-183] ^ d[511-180] ^ d[511-179] ^ d[511-169] ^ d[511-168] ^ d[511-167] ^ d[511-166] ^ d[511-164] ^ d[511-163] ^ d[511-159] ^ d[511-158] ^ d[511-155] ^ d[511-153] ^ d[511-152] ^ d[511-148] ^ d[511-146] ^ d[511-141] ^ d[511-140] ^ d[511-134] ^ d[511-133] ^ d[511-132] ^ d[511-131] ^ d[511-129] ^ d[511-125] ^ d[511-124] ^ d[511-123] ^ d[511-122] ^ d[511-120] ^ d[511-116] ^ d[511-115] ^ d[511-114] ^ d[511-113] ^ d[511-111] ^ d[511-110] ^ d[511-108] ^ d[511-107] ^ d[511-103] ^ d[511-101] ^ d[511-100] ^ d[511-98] ^ d[511-96] ^ d[511-95] ^ d[511-94] ^ d[511-93] ^ d[511-92] ^ d[511-91] ^ d[511-84] ^ d[511-82] ^ d[511-81] ^ d[511-80] ^ d[511-79] ^ d[511-78] ^ d[511-76] ^ d[511-70] ^ d[511-69] ^ d[511-65] ^ d[511-64] ^ d[511-63] ^ d[511-62] ^ d[511-60] ^ d[511-58] ^ d[511-57] ^ d[511-55] ^ d[511-52] ^ d[511-51] ^ d[511-50] ^ d[511-47] ^ d[511-45] ^ d[511-44] ^ d[511-42] ^ d[511-41] ^ d[511-34] ^ d[511-31] ^ d[511-29] ^ d[511-28] ^ d[511-27] ^ d[511-26] ^ d[511-25] ^ d[511-23] ^ d[511-22] ^ d[511-21] ^ d[511-13] ^ d[511-9] ^ d[511-7] ^ d[511-6] ^ d[511-3] ^ c[31-0] ^ c[31-3] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-17] ^ c[31-18] ^ c[31-19] ^ c[31-23] ^ c[31-24] ^ c[31-25] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-31];
                stage_crc512_crc[1] <= d[511-510] ^ d[511-509] ^ d[511-508] ^ d[511-506] ^ d[511-505] ^ d[511-504] ^ d[511-500] ^ d[511-499] ^ d[511-498] ^ d[511-493] ^ d[511-492] ^ d[511-491] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-487] ^ d[511-486] ^ d[511-484] ^ d[511-481] ^ d[511-480] ^ d[511-479] ^ d[511-478] ^ d[511-477] ^ d[511-475] ^ d[511-474] ^ d[511-470] ^ d[511-468] ^ d[511-466] ^ d[511-463] ^ d[511-462] ^ d[511-460] ^ d[511-459] ^ d[511-456] ^ d[511-450] ^ d[511-448] ^ d[511-447] ^ d[511-446] ^ d[511-442] ^ d[511-435] ^ d[511-434] ^ d[511-432] ^ d[511-431] ^ d[511-422] ^ d[511-420] ^ d[511-417] ^ d[511-416] ^ d[511-414] ^ d[511-412] ^ d[511-410] ^ d[511-407] ^ d[511-406] ^ d[511-405] ^ d[511-403] ^ d[511-402] ^ d[511-398] ^ d[511-397] ^ d[511-396] ^ d[511-394] ^ d[511-391] ^ d[511-390] ^ d[511-389] ^ d[511-388] ^ d[511-386] ^ d[511-385] ^ d[511-384] ^ d[511-379] ^ d[511-376] ^ d[511-374] ^ d[511-372] ^ d[511-370] ^ d[511-367] ^ d[511-366] ^ d[511-364] ^ d[511-361] ^ d[511-360] ^ d[511-357] ^ d[511-356] ^ d[511-355] ^ d[511-351] ^ d[511-347] ^ d[511-346] ^ d[511-345] ^ d[511-343] ^ d[511-342] ^ d[511-340] ^ d[511-339] ^ d[511-337] ^ d[511-336] ^ d[511-335] ^ d[511-333] ^ d[511-332] ^ d[511-331] ^ d[511-326] ^ d[511-325] ^ d[511-320] ^ d[511-319] ^ d[511-318] ^ d[511-317] ^ d[511-316] ^ d[511-315] ^ d[511-313] ^ d[511-310] ^ d[511-308] ^ d[511-307] ^ d[511-303] ^ d[511-301] ^ d[511-300] ^ d[511-298] ^ d[511-297] ^ d[511-296] ^ d[511-295] ^ d[511-294] ^ d[511-293] ^ d[511-292] ^ d[511-290] ^ d[511-288] ^ d[511-286] ^ d[511-285] ^ d[511-284] ^ d[511-281] ^ d[511-277] ^ d[511-275] ^ d[511-274] ^ d[511-272] ^ d[511-271] ^ d[511-267] ^ d[511-266] ^ d[511-263] ^ d[511-262] ^ d[511-259] ^ d[511-257] ^ d[511-255] ^ d[511-253] ^ d[511-250] ^ d[511-246] ^ d[511-241] ^ d[511-235] ^ d[511-232] ^ d[511-228] ^ d[511-226] ^ d[511-225] ^ d[511-224] ^ d[511-222] ^ d[511-214] ^ d[511-212] ^ d[511-210] ^ d[511-208] ^ d[511-207] ^ d[511-206] ^ d[511-205] ^ d[511-201] ^ d[511-200] ^ d[511-199] ^ d[511-197] ^ d[511-196] ^ d[511-195] ^ d[511-192] ^ d[511-191] ^ d[511-190] ^ d[511-189] ^ d[511-188] ^ d[511-186] ^ d[511-184] ^ d[511-181] ^ d[511-180] ^ d[511-170] ^ d[511-169] ^ d[511-168] ^ d[511-167] ^ d[511-165] ^ d[511-164] ^ d[511-160] ^ d[511-159] ^ d[511-156] ^ d[511-154] ^ d[511-153] ^ d[511-149] ^ d[511-147] ^ d[511-142] ^ d[511-141] ^ d[511-135] ^ d[511-134] ^ d[511-133] ^ d[511-132] ^ d[511-130] ^ d[511-126] ^ d[511-125] ^ d[511-124] ^ d[511-123] ^ d[511-121] ^ d[511-117] ^ d[511-116] ^ d[511-115] ^ d[511-114] ^ d[511-112] ^ d[511-111] ^ d[511-109] ^ d[511-108] ^ d[511-104] ^ d[511-102] ^ d[511-101] ^ d[511-99] ^ d[511-97] ^ d[511-96] ^ d[511-95] ^ d[511-94] ^ d[511-93] ^ d[511-92] ^ d[511-85] ^ d[511-83] ^ d[511-82] ^ d[511-81] ^ d[511-80] ^ d[511-79] ^ d[511-77] ^ d[511-71] ^ d[511-70] ^ d[511-66] ^ d[511-65] ^ d[511-64] ^ d[511-63] ^ d[511-61] ^ d[511-59] ^ d[511-58] ^ d[511-56] ^ d[511-53] ^ d[511-52] ^ d[511-51] ^ d[511-48] ^ d[511-46] ^ d[511-45] ^ d[511-43] ^ d[511-42] ^ d[511-35] ^ d[511-32] ^ d[511-30] ^ d[511-29] ^ d[511-28] ^ d[511-27] ^ d[511-26] ^ d[511-24] ^ d[511-23] ^ d[511-22] ^ d[511-14] ^ d[511-10] ^ d[511-8] ^ d[511-7] ^ d[511-4] ^ c[31-0] ^ c[31-1] ^ c[31-4] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-18] ^ c[31-19] ^ c[31-20] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-28] ^ c[31-29] ^ c[31-30];
                stage_crc512_crc[0] <= d[511-511] ^ d[511-510] ^ d[511-509] ^ d[511-507] ^ d[511-506] ^ d[511-505] ^ d[511-501] ^ d[511-500] ^ d[511-499] ^ d[511-494] ^ d[511-493] ^ d[511-492] ^ d[511-491] ^ d[511-490] ^ d[511-489] ^ d[511-488] ^ d[511-487] ^ d[511-485] ^ d[511-482] ^ d[511-481] ^ d[511-480] ^ d[511-479] ^ d[511-478] ^ d[511-476] ^ d[511-475] ^ d[511-471] ^ d[511-469] ^ d[511-467] ^ d[511-464] ^ d[511-463] ^ d[511-461] ^ d[511-460] ^ d[511-457] ^ d[511-451] ^ d[511-449] ^ d[511-448] ^ d[511-447] ^ d[511-443] ^ d[511-436] ^ d[511-435] ^ d[511-433] ^ d[511-432] ^ d[511-423] ^ d[511-421] ^ d[511-418] ^ d[511-417] ^ d[511-415] ^ d[511-413] ^ d[511-411] ^ d[511-408] ^ d[511-407] ^ d[511-406] ^ d[511-404] ^ d[511-403] ^ d[511-399] ^ d[511-398] ^ d[511-397] ^ d[511-395] ^ d[511-392] ^ d[511-391] ^ d[511-390] ^ d[511-389] ^ d[511-387] ^ d[511-386] ^ d[511-385] ^ d[511-380] ^ d[511-377] ^ d[511-375] ^ d[511-373] ^ d[511-371] ^ d[511-368] ^ d[511-367] ^ d[511-365] ^ d[511-362] ^ d[511-361] ^ d[511-358] ^ d[511-357] ^ d[511-356] ^ d[511-352] ^ d[511-348] ^ d[511-347] ^ d[511-346] ^ d[511-344] ^ d[511-343] ^ d[511-341] ^ d[511-340] ^ d[511-338] ^ d[511-337] ^ d[511-336] ^ d[511-334] ^ d[511-333] ^ d[511-332] ^ d[511-327] ^ d[511-326] ^ d[511-321] ^ d[511-320] ^ d[511-319] ^ d[511-318] ^ d[511-317] ^ d[511-316] ^ d[511-314] ^ d[511-311] ^ d[511-309] ^ d[511-308] ^ d[511-304] ^ d[511-302] ^ d[511-301] ^ d[511-299] ^ d[511-298] ^ d[511-297] ^ d[511-296] ^ d[511-295] ^ d[511-294] ^ d[511-293] ^ d[511-291] ^ d[511-289] ^ d[511-287] ^ d[511-286] ^ d[511-285] ^ d[511-282] ^ d[511-278] ^ d[511-276] ^ d[511-275] ^ d[511-273] ^ d[511-272] ^ d[511-268] ^ d[511-267] ^ d[511-264] ^ d[511-263] ^ d[511-260] ^ d[511-258] ^ d[511-256] ^ d[511-254] ^ d[511-251] ^ d[511-247] ^ d[511-242] ^ d[511-236] ^ d[511-233] ^ d[511-229] ^ d[511-227] ^ d[511-226] ^ d[511-225] ^ d[511-223] ^ d[511-215] ^ d[511-213] ^ d[511-211] ^ d[511-209] ^ d[511-208] ^ d[511-207] ^ d[511-206] ^ d[511-202] ^ d[511-201] ^ d[511-200] ^ d[511-198] ^ d[511-197] ^ d[511-196] ^ d[511-193] ^ d[511-192] ^ d[511-191] ^ d[511-190] ^ d[511-189] ^ d[511-187] ^ d[511-185] ^ d[511-182] ^ d[511-181] ^ d[511-171] ^ d[511-170] ^ d[511-169] ^ d[511-168] ^ d[511-166] ^ d[511-165] ^ d[511-161] ^ d[511-160] ^ d[511-157] ^ d[511-155] ^ d[511-154] ^ d[511-150] ^ d[511-148] ^ d[511-143] ^ d[511-142] ^ d[511-136] ^ d[511-135] ^ d[511-134] ^ d[511-133] ^ d[511-131] ^ d[511-127] ^ d[511-126] ^ d[511-125] ^ d[511-124] ^ d[511-122] ^ d[511-118] ^ d[511-117] ^ d[511-116] ^ d[511-115] ^ d[511-113] ^ d[511-112] ^ d[511-110] ^ d[511-109] ^ d[511-105] ^ d[511-103] ^ d[511-102] ^ d[511-100] ^ d[511-98] ^ d[511-97] ^ d[511-96] ^ d[511-95] ^ d[511-94] ^ d[511-93] ^ d[511-86] ^ d[511-84] ^ d[511-83] ^ d[511-82] ^ d[511-81] ^ d[511-80] ^ d[511-78] ^ d[511-72] ^ d[511-71] ^ d[511-67] ^ d[511-66] ^ d[511-65] ^ d[511-64] ^ d[511-62] ^ d[511-60] ^ d[511-59] ^ d[511-57] ^ d[511-54] ^ d[511-53] ^ d[511-52] ^ d[511-49] ^ d[511-47] ^ d[511-46] ^ d[511-44] ^ d[511-43] ^ d[511-36] ^ d[511-33] ^ d[511-31] ^ d[511-30] ^ d[511-29] ^ d[511-28] ^ d[511-27] ^ d[511-25] ^ d[511-24] ^ d[511-23] ^ d[511-15] ^ d[511-11] ^ d[511-9] ^ d[511-8] ^ d[511-5] ^ c[31-0] ^ c[31-1] ^ c[31-2] ^ c[31-5] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-19] ^ c[31-20] ^ c[31-21] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-29] ^ c[31-30] ^ c[31-31];

            end else if(stage_masking_keep == 64'h000000ffffffffff) begin

                // === CRC320 ===

                // Forward direct signals: valid, last, keep, data_bypass
                stage_crc320_valid <= stage_masking_valid; 
                stage_crc320_last <= stage_masking_last; 
                stage_crc320_keep <= stage_masking_keep; 
                stage_crc320_data_bypass <= stage_masking_data; 

                // Reset all other signals of the parallel CRC pipelines 
                stage_crc512_valid <= 1'b0; 
                stage_crc512_last <= 1'b0; 
                stage_crc512_keep <= 64'b0; 
                stage_crc512_data_bypass <= 512'b0; 
                stage_crc512_crc <= 32'b0; 

                for(integer pipeline_stage = 0; pipeline_stage < 16; pipeline_stage++) begin
                    stage_crc32_valid[pipeline_stage] <= 1'b0; 
                    stage_crc32_last[pipeline_stage] <= 1'b0; 
                    stage_crc32_keep[pipeline_stage] <= 64'b0; 
                    stage_crc32_data_bypass[pipeline_stage] <= 512'b0; 
                    stage_crc32_crc[pipeline_stage] <= 32'b0; 
                end 

                // Bitwise calculation of the CRC320-value based on the bitmasked data and the CRC-seed
                stage_crc320_crc[31] <= d[319-319] ^ d[319-318] ^ d[319-317] ^ d[319-315] ^ d[319-312] ^ d[319-310] ^ d[319-309] ^ d[319-305] ^ d[319-303] ^ d[319-302] ^ d[319-300] ^ d[319-299] ^ d[319-298] ^ d[319-297] ^ d[319-296] ^ d[319-295] ^ d[319-294] ^ d[319-292] ^ d[319-290] ^ d[319-288] ^ d[319-287] ^ d[319-286] ^ d[319-283] ^ d[319-279] ^ d[319-277] ^ d[319-276] ^ d[319-274] ^ d[319-273] ^ d[319-269] ^ d[319-268] ^ d[319-265] ^ d[319-264] ^ d[319-261] ^ d[319-259] ^ d[319-257] ^ d[319-255] ^ d[319-252] ^ d[319-248] ^ d[319-243] ^ d[319-237] ^ d[319-234] ^ d[319-230] ^ d[319-228] ^ d[319-227] ^ d[319-226] ^ d[319-224] ^ d[319-216] ^ d[319-214] ^ d[319-212] ^ d[319-210] ^ d[319-209] ^ d[319-208] ^ d[319-207] ^ d[319-203] ^ d[319-202] ^ d[319-201] ^ d[319-199] ^ d[319-198] ^ d[319-197] ^ d[319-194] ^ d[319-193] ^ d[319-192] ^ d[319-191] ^ d[319-190] ^ d[319-188] ^ d[319-186] ^ d[319-183] ^ d[319-182] ^ d[319-172] ^ d[319-171] ^ d[319-170] ^ d[319-169] ^ d[319-167] ^ d[319-166] ^ d[319-162] ^ d[319-161] ^ d[319-158] ^ d[319-156] ^ d[319-155] ^ d[319-151] ^ d[319-149] ^ d[319-144] ^ d[319-143] ^ d[319-137] ^ d[319-136] ^ d[319-135] ^ d[319-134] ^ d[319-132] ^ d[319-128] ^ d[319-127] ^ d[319-126] ^ d[319-125] ^ d[319-123] ^ d[319-119] ^ d[319-118] ^ d[319-117] ^ d[319-116] ^ d[319-114] ^ d[319-113] ^ d[319-111] ^ d[319-110] ^ d[319-106] ^ d[319-104] ^ d[319-103] ^ d[319-101] ^ d[319-99] ^ d[319-98] ^ d[319-97] ^ d[319-96] ^ d[319-95] ^ d[319-94] ^ d[319-87] ^ d[319-85] ^ d[319-84] ^ d[319-83] ^ d[319-82] ^ d[319-81] ^ d[319-79] ^ d[319-73] ^ d[319-72] ^ d[319-68] ^ d[319-67] ^ d[319-66] ^ d[319-65] ^ d[319-63] ^ d[319-61] ^ d[319-60] ^ d[319-58] ^ d[319-55] ^ d[319-54] ^ d[319-53] ^ d[319-50] ^ d[319-48] ^ d[319-47] ^ d[319-45] ^ d[319-44] ^ d[319-37] ^ d[319-34] ^ d[319-32] ^ d[319-31] ^ d[319-30] ^ d[319-29] ^ d[319-28] ^ d[319-26] ^ d[319-25] ^ d[319-24] ^ d[319-16] ^ d[319-12] ^ d[319-10] ^ d[319-9] ^ d[319-6] ^ d[319-0] ^ c[31-0] ^ c[31-2] ^ c[31-4] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-14] ^ c[31-15] ^ c[31-17] ^ c[31-21] ^ c[31-22] ^ c[31-24] ^ c[31-27] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc320_crc[30] <= d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-313] ^ d[319-312] ^ d[319-311] ^ d[319-309] ^ d[319-306] ^ d[319-305] ^ d[319-304] ^ d[319-302] ^ d[319-301] ^ d[319-294] ^ d[319-293] ^ d[319-292] ^ d[319-291] ^ d[319-290] ^ d[319-289] ^ d[319-286] ^ d[319-284] ^ d[319-283] ^ d[319-280] ^ d[319-279] ^ d[319-278] ^ d[319-276] ^ d[319-275] ^ d[319-273] ^ d[319-270] ^ d[319-268] ^ d[319-266] ^ d[319-264] ^ d[319-262] ^ d[319-261] ^ d[319-260] ^ d[319-259] ^ d[319-258] ^ d[319-257] ^ d[319-256] ^ d[319-255] ^ d[319-253] ^ d[319-252] ^ d[319-249] ^ d[319-248] ^ d[319-244] ^ d[319-243] ^ d[319-238] ^ d[319-237] ^ d[319-235] ^ d[319-234] ^ d[319-231] ^ d[319-230] ^ d[319-229] ^ d[319-226] ^ d[319-225] ^ d[319-224] ^ d[319-217] ^ d[319-216] ^ d[319-215] ^ d[319-214] ^ d[319-213] ^ d[319-212] ^ d[319-211] ^ d[319-207] ^ d[319-204] ^ d[319-201] ^ d[319-200] ^ d[319-197] ^ d[319-195] ^ d[319-190] ^ d[319-189] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-184] ^ d[319-182] ^ d[319-173] ^ d[319-169] ^ d[319-168] ^ d[319-166] ^ d[319-163] ^ d[319-161] ^ d[319-159] ^ d[319-158] ^ d[319-157] ^ d[319-155] ^ d[319-152] ^ d[319-151] ^ d[319-150] ^ d[319-149] ^ d[319-145] ^ d[319-143] ^ d[319-138] ^ d[319-134] ^ d[319-133] ^ d[319-132] ^ d[319-129] ^ d[319-125] ^ d[319-124] ^ d[319-123] ^ d[319-120] ^ d[319-116] ^ d[319-115] ^ d[319-113] ^ d[319-112] ^ d[319-110] ^ d[319-107] ^ d[319-106] ^ d[319-105] ^ d[319-103] ^ d[319-102] ^ d[319-101] ^ d[319-100] ^ d[319-94] ^ d[319-88] ^ d[319-87] ^ d[319-86] ^ d[319-81] ^ d[319-80] ^ d[319-79] ^ d[319-74] ^ d[319-72] ^ d[319-69] ^ d[319-65] ^ d[319-64] ^ d[319-63] ^ d[319-62] ^ d[319-60] ^ d[319-59] ^ d[319-58] ^ d[319-56] ^ d[319-53] ^ d[319-51] ^ d[319-50] ^ d[319-49] ^ d[319-47] ^ d[319-46] ^ d[319-44] ^ d[319-38] ^ d[319-37] ^ d[319-35] ^ d[319-34] ^ d[319-33] ^ d[319-28] ^ d[319-27] ^ d[319-24] ^ d[319-17] ^ d[319-16] ^ d[319-13] ^ d[319-12] ^ d[319-11] ^ d[319-9] ^ d[319-7] ^ d[319-6] ^ d[319-1] ^ d[319-0] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-13] ^ c[31-14] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-21] ^ c[31-23] ^ c[31-24] ^ c[31-25] ^ c[31-27] ^ c[31-28] ^ c[31-29];
                stage_crc320_crc[29] <= d[319-319] ^ d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-313] ^ d[319-309] ^ d[319-307] ^ d[319-306] ^ d[319-300] ^ d[319-299] ^ d[319-298] ^ d[319-297] ^ d[319-296] ^ d[319-293] ^ d[319-291] ^ d[319-288] ^ d[319-286] ^ d[319-285] ^ d[319-284] ^ d[319-283] ^ d[319-281] ^ d[319-280] ^ d[319-273] ^ d[319-271] ^ d[319-268] ^ d[319-267] ^ d[319-264] ^ d[319-263] ^ d[319-262] ^ d[319-260] ^ d[319-258] ^ d[319-256] ^ d[319-255] ^ d[319-254] ^ d[319-253] ^ d[319-252] ^ d[319-250] ^ d[319-249] ^ d[319-248] ^ d[319-245] ^ d[319-244] ^ d[319-243] ^ d[319-239] ^ d[319-238] ^ d[319-237] ^ d[319-236] ^ d[319-235] ^ d[319-234] ^ d[319-232] ^ d[319-231] ^ d[319-228] ^ d[319-225] ^ d[319-224] ^ d[319-218] ^ d[319-217] ^ d[319-215] ^ d[319-213] ^ d[319-210] ^ d[319-209] ^ d[319-207] ^ d[319-205] ^ d[319-203] ^ d[319-199] ^ d[319-197] ^ d[319-196] ^ d[319-194] ^ d[319-193] ^ d[319-192] ^ d[319-189] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-182] ^ d[319-174] ^ d[319-172] ^ d[319-171] ^ d[319-166] ^ d[319-164] ^ d[319-161] ^ d[319-160] ^ d[319-159] ^ d[319-155] ^ d[319-153] ^ d[319-152] ^ d[319-150] ^ d[319-149] ^ d[319-146] ^ d[319-143] ^ d[319-139] ^ d[319-137] ^ d[319-136] ^ d[319-133] ^ d[319-132] ^ d[319-130] ^ d[319-128] ^ d[319-127] ^ d[319-124] ^ d[319-123] ^ d[319-121] ^ d[319-119] ^ d[319-118] ^ d[319-110] ^ d[319-108] ^ d[319-107] ^ d[319-102] ^ d[319-99] ^ d[319-98] ^ d[319-97] ^ d[319-96] ^ d[319-94] ^ d[319-89] ^ d[319-88] ^ d[319-85] ^ d[319-84] ^ d[319-83] ^ d[319-80] ^ d[319-79] ^ d[319-75] ^ d[319-72] ^ d[319-70] ^ d[319-68] ^ d[319-67] ^ d[319-64] ^ d[319-59] ^ d[319-58] ^ d[319-57] ^ d[319-55] ^ d[319-53] ^ d[319-52] ^ d[319-51] ^ d[319-44] ^ d[319-39] ^ d[319-38] ^ d[319-37] ^ d[319-36] ^ d[319-35] ^ d[319-32] ^ d[319-31] ^ d[319-30] ^ d[319-26] ^ d[319-24] ^ d[319-18] ^ d[319-17] ^ d[319-16] ^ d[319-14] ^ d[319-13] ^ d[319-9] ^ d[319-8] ^ d[319-7] ^ d[319-6] ^ d[319-2] ^ d[319-1] ^ d[319-0] ^ c[31-0] ^ c[31-3] ^ c[31-5] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-18] ^ c[31-19] ^ c[31-21] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-31];
                stage_crc320_crc[28] <= d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-310] ^ d[319-308] ^ d[319-307] ^ d[319-301] ^ d[319-300] ^ d[319-299] ^ d[319-298] ^ d[319-297] ^ d[319-294] ^ d[319-292] ^ d[319-289] ^ d[319-287] ^ d[319-286] ^ d[319-285] ^ d[319-284] ^ d[319-282] ^ d[319-281] ^ d[319-274] ^ d[319-272] ^ d[319-269] ^ d[319-268] ^ d[319-265] ^ d[319-264] ^ d[319-263] ^ d[319-261] ^ d[319-259] ^ d[319-257] ^ d[319-256] ^ d[319-255] ^ d[319-254] ^ d[319-253] ^ d[319-251] ^ d[319-250] ^ d[319-249] ^ d[319-246] ^ d[319-245] ^ d[319-244] ^ d[319-240] ^ d[319-239] ^ d[319-238] ^ d[319-237] ^ d[319-236] ^ d[319-235] ^ d[319-233] ^ d[319-232] ^ d[319-229] ^ d[319-226] ^ d[319-225] ^ d[319-219] ^ d[319-218] ^ d[319-216] ^ d[319-214] ^ d[319-211] ^ d[319-210] ^ d[319-208] ^ d[319-206] ^ d[319-204] ^ d[319-200] ^ d[319-198] ^ d[319-197] ^ d[319-195] ^ d[319-194] ^ d[319-193] ^ d[319-190] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-183] ^ d[319-175] ^ d[319-173] ^ d[319-172] ^ d[319-167] ^ d[319-165] ^ d[319-162] ^ d[319-161] ^ d[319-160] ^ d[319-156] ^ d[319-154] ^ d[319-153] ^ d[319-151] ^ d[319-150] ^ d[319-147] ^ d[319-144] ^ d[319-140] ^ d[319-138] ^ d[319-137] ^ d[319-134] ^ d[319-133] ^ d[319-131] ^ d[319-129] ^ d[319-128] ^ d[319-125] ^ d[319-124] ^ d[319-122] ^ d[319-120] ^ d[319-119] ^ d[319-111] ^ d[319-109] ^ d[319-108] ^ d[319-103] ^ d[319-100] ^ d[319-99] ^ d[319-98] ^ d[319-97] ^ d[319-95] ^ d[319-90] ^ d[319-89] ^ d[319-86] ^ d[319-85] ^ d[319-84] ^ d[319-81] ^ d[319-80] ^ d[319-76] ^ d[319-73] ^ d[319-71] ^ d[319-69] ^ d[319-68] ^ d[319-65] ^ d[319-60] ^ d[319-59] ^ d[319-58] ^ d[319-56] ^ d[319-54] ^ d[319-53] ^ d[319-52] ^ d[319-45] ^ d[319-40] ^ d[319-39] ^ d[319-38] ^ d[319-37] ^ d[319-36] ^ d[319-33] ^ d[319-32] ^ d[319-31] ^ d[319-27] ^ d[319-25] ^ d[319-19] ^ d[319-18] ^ d[319-17] ^ d[319-15] ^ d[319-14] ^ d[319-10] ^ d[319-9] ^ d[319-8] ^ d[319-7] ^ d[319-3] ^ d[319-2] ^ d[319-1] ^ c[31-1] ^ c[31-4] ^ c[31-6] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-19] ^ c[31-20] ^ c[31-22] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29];
                stage_crc320_crc[27] <= d[319-319] ^ d[319-316] ^ d[319-312] ^ d[319-311] ^ d[319-310] ^ d[319-308] ^ d[319-305] ^ d[319-303] ^ d[319-301] ^ d[319-297] ^ d[319-296] ^ d[319-294] ^ d[319-293] ^ d[319-292] ^ d[319-285] ^ d[319-282] ^ d[319-279] ^ d[319-277] ^ d[319-276] ^ d[319-275] ^ d[319-274] ^ d[319-270] ^ d[319-268] ^ d[319-266] ^ d[319-262] ^ d[319-261] ^ d[319-260] ^ d[319-259] ^ d[319-258] ^ d[319-256] ^ d[319-254] ^ d[319-251] ^ d[319-250] ^ d[319-248] ^ d[319-247] ^ d[319-246] ^ d[319-245] ^ d[319-243] ^ d[319-241] ^ d[319-240] ^ d[319-239] ^ d[319-238] ^ d[319-236] ^ d[319-233] ^ d[319-228] ^ d[319-224] ^ d[319-220] ^ d[319-219] ^ d[319-217] ^ d[319-216] ^ d[319-215] ^ d[319-214] ^ d[319-211] ^ d[319-210] ^ d[319-208] ^ d[319-205] ^ d[319-203] ^ d[319-202] ^ d[319-197] ^ d[319-196] ^ d[319-195] ^ d[319-193] ^ d[319-192] ^ d[319-190] ^ d[319-189] ^ d[319-187] ^ d[319-186] ^ d[319-184] ^ d[319-183] ^ d[319-182] ^ d[319-176] ^ d[319-174] ^ d[319-173] ^ d[319-172] ^ d[319-171] ^ d[319-170] ^ d[319-169] ^ d[319-168] ^ d[319-167] ^ d[319-163] ^ d[319-158] ^ d[319-157] ^ d[319-156] ^ d[319-154] ^ d[319-152] ^ d[319-149] ^ d[319-148] ^ d[319-145] ^ d[319-144] ^ d[319-143] ^ d[319-141] ^ d[319-139] ^ d[319-138] ^ d[319-137] ^ d[319-136] ^ d[319-130] ^ d[319-129] ^ d[319-128] ^ d[319-127] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-118] ^ d[319-117] ^ d[319-116] ^ d[319-114] ^ d[319-113] ^ d[319-112] ^ d[319-111] ^ d[319-109] ^ d[319-106] ^ d[319-103] ^ d[319-100] ^ d[319-97] ^ d[319-95] ^ d[319-94] ^ d[319-91] ^ d[319-90] ^ d[319-86] ^ d[319-84] ^ d[319-83] ^ d[319-79] ^ d[319-77] ^ d[319-74] ^ d[319-73] ^ d[319-70] ^ d[319-69] ^ d[319-68] ^ d[319-67] ^ d[319-65] ^ d[319-63] ^ d[319-59] ^ d[319-58] ^ d[319-57] ^ d[319-50] ^ d[319-48] ^ d[319-47] ^ d[319-46] ^ d[319-45] ^ d[319-44] ^ d[319-41] ^ d[319-40] ^ d[319-39] ^ d[319-38] ^ d[319-33] ^ d[319-31] ^ d[319-30] ^ d[319-29] ^ d[319-25] ^ d[319-24] ^ d[319-20] ^ d[319-19] ^ d[319-18] ^ d[319-15] ^ d[319-12] ^ d[319-11] ^ d[319-8] ^ d[319-6] ^ d[319-4] ^ d[319-3] ^ d[319-2] ^ d[319-0] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-8] ^ c[31-9] ^ c[31-13] ^ c[31-15] ^ c[31-17] ^ c[31-20] ^ c[31-22] ^ c[31-23] ^ c[31-24] ^ c[31-28] ^ c[31-31];
                stage_crc320_crc[26] <= d[319-319] ^ d[319-318] ^ d[319-315] ^ d[319-313] ^ d[319-311] ^ d[319-310] ^ d[319-306] ^ d[319-305] ^ d[319-304] ^ d[319-303] ^ d[319-300] ^ d[319-299] ^ d[319-296] ^ d[319-293] ^ d[319-292] ^ d[319-290] ^ d[319-288] ^ d[319-287] ^ d[319-280] ^ d[319-279] ^ d[319-278] ^ d[319-275] ^ d[319-274] ^ d[319-273] ^ d[319-271] ^ d[319-268] ^ d[319-267] ^ d[319-265] ^ d[319-264] ^ d[319-263] ^ d[319-262] ^ d[319-260] ^ d[319-251] ^ d[319-249] ^ d[319-247] ^ d[319-246] ^ d[319-244] ^ d[319-243] ^ d[319-242] ^ d[319-241] ^ d[319-240] ^ d[319-239] ^ d[319-230] ^ d[319-229] ^ d[319-228] ^ d[319-227] ^ d[319-226] ^ d[319-225] ^ d[319-224] ^ d[319-221] ^ d[319-220] ^ d[319-218] ^ d[319-217] ^ d[319-215] ^ d[319-214] ^ d[319-211] ^ d[319-210] ^ d[319-208] ^ d[319-207] ^ d[319-206] ^ d[319-204] ^ d[319-202] ^ d[319-201] ^ d[319-199] ^ d[319-196] ^ d[319-192] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-184] ^ d[319-182] ^ d[319-177] ^ d[319-175] ^ d[319-174] ^ d[319-173] ^ d[319-168] ^ d[319-167] ^ d[319-166] ^ d[319-164] ^ d[319-162] ^ d[319-161] ^ d[319-159] ^ d[319-157] ^ d[319-156] ^ d[319-153] ^ d[319-151] ^ d[319-150] ^ d[319-146] ^ d[319-145] ^ d[319-143] ^ d[319-142] ^ d[319-140] ^ d[319-139] ^ d[319-138] ^ d[319-136] ^ d[319-135] ^ d[319-134] ^ d[319-132] ^ d[319-131] ^ d[319-130] ^ d[319-129] ^ d[319-127] ^ d[319-126] ^ d[319-125] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-116] ^ d[319-115] ^ d[319-112] ^ d[319-111] ^ d[319-107] ^ d[319-106] ^ d[319-103] ^ d[319-99] ^ d[319-97] ^ d[319-94] ^ d[319-92] ^ d[319-91] ^ d[319-83] ^ d[319-82] ^ d[319-81] ^ d[319-80] ^ d[319-79] ^ d[319-78] ^ d[319-75] ^ d[319-74] ^ d[319-73] ^ d[319-72] ^ d[319-71] ^ d[319-70] ^ d[319-69] ^ d[319-67] ^ d[319-65] ^ d[319-64] ^ d[319-63] ^ d[319-61] ^ d[319-59] ^ d[319-55] ^ d[319-54] ^ d[319-53] ^ d[319-51] ^ d[319-50] ^ d[319-49] ^ d[319-46] ^ d[319-44] ^ d[319-42] ^ d[319-41] ^ d[319-40] ^ d[319-39] ^ d[319-37] ^ d[319-29] ^ d[319-28] ^ d[319-24] ^ d[319-21] ^ d[319-20] ^ d[319-19] ^ d[319-13] ^ d[319-10] ^ d[319-7] ^ d[319-6] ^ d[319-5] ^ d[319-4] ^ d[319-3] ^ d[319-1] ^ d[319-0] ^ c[31-0] ^ c[31-2] ^ c[31-4] ^ c[31-5] ^ c[31-8] ^ c[31-11] ^ c[31-12] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-22] ^ c[31-23] ^ c[31-25] ^ c[31-27] ^ c[31-30] ^ c[31-31];
                stage_crc320_crc[25] <= d[319-319] ^ d[319-316] ^ d[319-314] ^ d[319-312] ^ d[319-311] ^ d[319-307] ^ d[319-306] ^ d[319-305] ^ d[319-304] ^ d[319-301] ^ d[319-300] ^ d[319-297] ^ d[319-294] ^ d[319-293] ^ d[319-291] ^ d[319-289] ^ d[319-288] ^ d[319-281] ^ d[319-280] ^ d[319-279] ^ d[319-276] ^ d[319-275] ^ d[319-274] ^ d[319-272] ^ d[319-269] ^ d[319-268] ^ d[319-266] ^ d[319-265] ^ d[319-264] ^ d[319-263] ^ d[319-261] ^ d[319-252] ^ d[319-250] ^ d[319-248] ^ d[319-247] ^ d[319-245] ^ d[319-244] ^ d[319-243] ^ d[319-242] ^ d[319-241] ^ d[319-240] ^ d[319-231] ^ d[319-230] ^ d[319-229] ^ d[319-228] ^ d[319-227] ^ d[319-226] ^ d[319-225] ^ d[319-222] ^ d[319-221] ^ d[319-219] ^ d[319-218] ^ d[319-216] ^ d[319-215] ^ d[319-212] ^ d[319-211] ^ d[319-209] ^ d[319-208] ^ d[319-207] ^ d[319-205] ^ d[319-203] ^ d[319-202] ^ d[319-200] ^ d[319-197] ^ d[319-193] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-183] ^ d[319-178] ^ d[319-176] ^ d[319-175] ^ d[319-174] ^ d[319-169] ^ d[319-168] ^ d[319-167] ^ d[319-165] ^ d[319-163] ^ d[319-162] ^ d[319-160] ^ d[319-158] ^ d[319-157] ^ d[319-154] ^ d[319-152] ^ d[319-151] ^ d[319-147] ^ d[319-146] ^ d[319-144] ^ d[319-143] ^ d[319-141] ^ d[319-140] ^ d[319-139] ^ d[319-137] ^ d[319-136] ^ d[319-135] ^ d[319-133] ^ d[319-132] ^ d[319-131] ^ d[319-130] ^ d[319-128] ^ d[319-127] ^ d[319-126] ^ d[319-124] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-117] ^ d[319-116] ^ d[319-113] ^ d[319-112] ^ d[319-108] ^ d[319-107] ^ d[319-104] ^ d[319-100] ^ d[319-98] ^ d[319-95] ^ d[319-93] ^ d[319-92] ^ d[319-84] ^ d[319-83] ^ d[319-82] ^ d[319-81] ^ d[319-80] ^ d[319-79] ^ d[319-76] ^ d[319-75] ^ d[319-74] ^ d[319-73] ^ d[319-72] ^ d[319-71] ^ d[319-70] ^ d[319-68] ^ d[319-66] ^ d[319-65] ^ d[319-64] ^ d[319-62] ^ d[319-60] ^ d[319-56] ^ d[319-55] ^ d[319-54] ^ d[319-52] ^ d[319-51] ^ d[319-50] ^ d[319-47] ^ d[319-45] ^ d[319-43] ^ d[319-42] ^ d[319-41] ^ d[319-40] ^ d[319-38] ^ d[319-30] ^ d[319-29] ^ d[319-25] ^ d[319-22] ^ d[319-21] ^ d[319-20] ^ d[319-14] ^ d[319-11] ^ d[319-8] ^ d[319-7] ^ d[319-6] ^ d[319-5] ^ d[319-4] ^ d[319-2] ^ d[319-1] ^ c[31-0] ^ c[31-1] ^ c[31-3] ^ c[31-5] ^ c[31-6] ^ c[31-9] ^ c[31-12] ^ c[31-13] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-19] ^ c[31-23] ^ c[31-24] ^ c[31-26] ^ c[31-28] ^ c[31-31];
                stage_crc320_crc[24] <= d[319-319] ^ d[319-318] ^ d[319-313] ^ d[319-310] ^ d[319-309] ^ d[319-308] ^ d[319-307] ^ d[319-306] ^ d[319-303] ^ d[319-301] ^ d[319-300] ^ d[319-299] ^ d[319-297] ^ d[319-296] ^ d[319-289] ^ d[319-288] ^ d[319-287] ^ d[319-286] ^ d[319-283] ^ d[319-282] ^ d[319-281] ^ d[319-280] ^ d[319-279] ^ d[319-275] ^ d[319-274] ^ d[319-270] ^ d[319-268] ^ d[319-267] ^ d[319-266] ^ d[319-262] ^ d[319-261] ^ d[319-259] ^ d[319-257] ^ d[319-255] ^ d[319-253] ^ d[319-252] ^ d[319-251] ^ d[319-249] ^ d[319-246] ^ d[319-245] ^ d[319-244] ^ d[319-242] ^ d[319-241] ^ d[319-237] ^ d[319-234] ^ d[319-232] ^ d[319-231] ^ d[319-229] ^ d[319-224] ^ d[319-223] ^ d[319-222] ^ d[319-220] ^ d[319-219] ^ d[319-217] ^ d[319-214] ^ d[319-213] ^ d[319-207] ^ d[319-206] ^ d[319-204] ^ d[319-202] ^ d[319-199] ^ d[319-197] ^ d[319-193] ^ d[319-192] ^ d[319-191] ^ d[319-190] ^ d[319-189] ^ d[319-187] ^ d[319-184] ^ d[319-183] ^ d[319-182] ^ d[319-179] ^ d[319-177] ^ d[319-176] ^ d[319-175] ^ d[319-172] ^ d[319-171] ^ d[319-168] ^ d[319-167] ^ d[319-164] ^ d[319-163] ^ d[319-162] ^ d[319-159] ^ d[319-156] ^ d[319-153] ^ d[319-152] ^ d[319-151] ^ d[319-149] ^ d[319-148] ^ d[319-147] ^ d[319-145] ^ d[319-143] ^ d[319-142] ^ d[319-141] ^ d[319-140] ^ d[319-138] ^ d[319-135] ^ d[319-133] ^ d[319-131] ^ d[319-129] ^ d[319-126] ^ d[319-124] ^ d[319-122] ^ d[319-119] ^ d[319-116] ^ d[319-111] ^ d[319-110] ^ d[319-109] ^ d[319-108] ^ d[319-106] ^ d[319-105] ^ d[319-104] ^ d[319-103] ^ d[319-98] ^ d[319-97] ^ d[319-95] ^ d[319-93] ^ d[319-87] ^ d[319-80] ^ d[319-79] ^ d[319-77] ^ d[319-76] ^ d[319-75] ^ d[319-74] ^ d[319-71] ^ d[319-69] ^ d[319-68] ^ d[319-60] ^ d[319-58] ^ d[319-57] ^ d[319-56] ^ d[319-54] ^ d[319-52] ^ d[319-51] ^ d[319-50] ^ d[319-47] ^ d[319-46] ^ d[319-45] ^ d[319-43] ^ d[319-42] ^ d[319-41] ^ d[319-39] ^ d[319-37] ^ d[319-34] ^ d[319-32] ^ d[319-29] ^ d[319-28] ^ d[319-25] ^ d[319-24] ^ d[319-23] ^ d[319-22] ^ d[319-21] ^ d[319-16] ^ d[319-15] ^ d[319-10] ^ d[319-8] ^ d[319-7] ^ d[319-5] ^ d[319-3] ^ d[319-2] ^ d[319-0] ^ c[31-0] ^ c[31-1] ^ c[31-8] ^ c[31-9] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-15] ^ c[31-18] ^ c[31-19] ^ c[31-20] ^ c[31-21] ^ c[31-22] ^ c[31-25] ^ c[31-30] ^ c[31-31];
                stage_crc320_crc[23] <= d[319-318] ^ d[319-317] ^ d[319-315] ^ d[319-314] ^ d[319-312] ^ d[319-311] ^ d[319-308] ^ d[319-307] ^ d[319-305] ^ d[319-304] ^ d[319-303] ^ d[319-301] ^ d[319-299] ^ d[319-296] ^ d[319-295] ^ d[319-294] ^ d[319-292] ^ d[319-289] ^ d[319-286] ^ d[319-284] ^ d[319-282] ^ d[319-281] ^ d[319-280] ^ d[319-279] ^ d[319-277] ^ d[319-275] ^ d[319-274] ^ d[319-273] ^ d[319-271] ^ d[319-267] ^ d[319-265] ^ d[319-264] ^ d[319-263] ^ d[319-262] ^ d[319-261] ^ d[319-260] ^ d[319-259] ^ d[319-258] ^ d[319-257] ^ d[319-256] ^ d[319-255] ^ d[319-254] ^ d[319-253] ^ d[319-250] ^ d[319-248] ^ d[319-247] ^ d[319-246] ^ d[319-245] ^ d[319-242] ^ d[319-238] ^ d[319-237] ^ d[319-235] ^ d[319-234] ^ d[319-233] ^ d[319-232] ^ d[319-228] ^ d[319-227] ^ d[319-226] ^ d[319-225] ^ d[319-223] ^ d[319-221] ^ d[319-220] ^ d[319-218] ^ d[319-216] ^ d[319-215] ^ d[319-212] ^ d[319-210] ^ d[319-209] ^ d[319-205] ^ d[319-202] ^ d[319-201] ^ d[319-200] ^ d[319-199] ^ d[319-197] ^ d[319-186] ^ d[319-185] ^ d[319-184] ^ d[319-182] ^ d[319-180] ^ d[319-178] ^ d[319-177] ^ d[319-176] ^ d[319-173] ^ d[319-171] ^ d[319-170] ^ d[319-168] ^ d[319-167] ^ d[319-166] ^ d[319-165] ^ d[319-164] ^ d[319-163] ^ d[319-162] ^ d[319-161] ^ d[319-160] ^ d[319-158] ^ d[319-157] ^ d[319-156] ^ d[319-155] ^ d[319-154] ^ d[319-153] ^ d[319-152] ^ d[319-151] ^ d[319-150] ^ d[319-148] ^ d[319-146] ^ d[319-142] ^ d[319-141] ^ d[319-139] ^ d[319-137] ^ d[319-135] ^ d[319-130] ^ d[319-128] ^ d[319-126] ^ d[319-120] ^ d[319-119] ^ d[319-118] ^ d[319-116] ^ d[319-114] ^ d[319-113] ^ d[319-112] ^ d[319-109] ^ d[319-107] ^ d[319-105] ^ d[319-103] ^ d[319-101] ^ d[319-97] ^ d[319-95] ^ d[319-88] ^ d[319-87] ^ d[319-85] ^ d[319-84] ^ d[319-83] ^ d[319-82] ^ d[319-80] ^ d[319-79] ^ d[319-78] ^ d[319-77] ^ d[319-76] ^ d[319-75] ^ d[319-73] ^ d[319-70] ^ d[319-69] ^ d[319-68] ^ d[319-67] ^ d[319-66] ^ d[319-65] ^ d[319-63] ^ d[319-60] ^ d[319-59] ^ d[319-57] ^ d[319-54] ^ d[319-52] ^ d[319-51] ^ d[319-50] ^ d[319-46] ^ d[319-45] ^ d[319-43] ^ d[319-42] ^ d[319-40] ^ d[319-38] ^ d[319-37] ^ d[319-35] ^ d[319-34] ^ d[319-33] ^ d[319-32] ^ d[319-31] ^ d[319-28] ^ d[319-23] ^ d[319-22] ^ d[319-17] ^ d[319-12] ^ d[319-11] ^ d[319-10] ^ d[319-8] ^ d[319-4] ^ d[319-3] ^ d[319-1] ^ d[319-0] ^ c[31-1] ^ c[31-4] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-11] ^ c[31-13] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-19] ^ c[31-20] ^ c[31-23] ^ c[31-24] ^ c[31-26] ^ c[31-27] ^ c[31-29] ^ c[31-30];
                stage_crc320_crc[22] <= d[319-319] ^ d[319-318] ^ d[319-316] ^ d[319-315] ^ d[319-313] ^ d[319-312] ^ d[319-309] ^ d[319-308] ^ d[319-306] ^ d[319-305] ^ d[319-304] ^ d[319-302] ^ d[319-300] ^ d[319-297] ^ d[319-296] ^ d[319-295] ^ d[319-293] ^ d[319-290] ^ d[319-287] ^ d[319-285] ^ d[319-283] ^ d[319-282] ^ d[319-281] ^ d[319-280] ^ d[319-278] ^ d[319-276] ^ d[319-275] ^ d[319-274] ^ d[319-272] ^ d[319-268] ^ d[319-266] ^ d[319-265] ^ d[319-264] ^ d[319-263] ^ d[319-262] ^ d[319-261] ^ d[319-260] ^ d[319-259] ^ d[319-258] ^ d[319-257] ^ d[319-256] ^ d[319-255] ^ d[319-254] ^ d[319-251] ^ d[319-249] ^ d[319-248] ^ d[319-247] ^ d[319-246] ^ d[319-243] ^ d[319-239] ^ d[319-238] ^ d[319-236] ^ d[319-235] ^ d[319-234] ^ d[319-233] ^ d[319-229] ^ d[319-228] ^ d[319-227] ^ d[319-226] ^ d[319-224] ^ d[319-222] ^ d[319-221] ^ d[319-219] ^ d[319-217] ^ d[319-216] ^ d[319-213] ^ d[319-211] ^ d[319-210] ^ d[319-206] ^ d[319-203] ^ d[319-202] ^ d[319-201] ^ d[319-200] ^ d[319-198] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-183] ^ d[319-181] ^ d[319-179] ^ d[319-178] ^ d[319-177] ^ d[319-174] ^ d[319-172] ^ d[319-171] ^ d[319-169] ^ d[319-168] ^ d[319-167] ^ d[319-166] ^ d[319-165] ^ d[319-164] ^ d[319-163] ^ d[319-162] ^ d[319-161] ^ d[319-159] ^ d[319-158] ^ d[319-157] ^ d[319-156] ^ d[319-155] ^ d[319-154] ^ d[319-153] ^ d[319-152] ^ d[319-151] ^ d[319-149] ^ d[319-147] ^ d[319-143] ^ d[319-142] ^ d[319-140] ^ d[319-138] ^ d[319-136] ^ d[319-131] ^ d[319-129] ^ d[319-127] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-117] ^ d[319-115] ^ d[319-114] ^ d[319-113] ^ d[319-110] ^ d[319-108] ^ d[319-106] ^ d[319-104] ^ d[319-102] ^ d[319-98] ^ d[319-96] ^ d[319-89] ^ d[319-88] ^ d[319-86] ^ d[319-85] ^ d[319-84] ^ d[319-83] ^ d[319-81] ^ d[319-80] ^ d[319-79] ^ d[319-78] ^ d[319-77] ^ d[319-76] ^ d[319-74] ^ d[319-71] ^ d[319-70] ^ d[319-69] ^ d[319-68] ^ d[319-67] ^ d[319-66] ^ d[319-64] ^ d[319-61] ^ d[319-60] ^ d[319-58] ^ d[319-55] ^ d[319-53] ^ d[319-52] ^ d[319-51] ^ d[319-47] ^ d[319-46] ^ d[319-44] ^ d[319-43] ^ d[319-41] ^ d[319-39] ^ d[319-38] ^ d[319-36] ^ d[319-35] ^ d[319-34] ^ d[319-33] ^ d[319-32] ^ d[319-29] ^ d[319-24] ^ d[319-23] ^ d[319-18] ^ d[319-13] ^ d[319-12] ^ d[319-11] ^ d[319-9] ^ d[319-5] ^ d[319-4] ^ d[319-2] ^ d[319-1] ^ c[31-2] ^ c[31-5] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-12] ^ c[31-14] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-20] ^ c[31-21] ^ c[31-24] ^ c[31-25] ^ c[31-27] ^ c[31-28] ^ c[31-30] ^ c[31-31];
                stage_crc320_crc[21] <= d[319-318] ^ d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-313] ^ d[319-312] ^ d[319-307] ^ d[319-306] ^ d[319-302] ^ d[319-301] ^ d[319-300] ^ d[319-299] ^ d[319-295] ^ d[319-292] ^ d[319-291] ^ d[319-290] ^ d[319-287] ^ d[319-284] ^ d[319-282] ^ d[319-281] ^ d[319-275] ^ d[319-274] ^ d[319-268] ^ d[319-267] ^ d[319-266] ^ d[319-263] ^ d[319-262] ^ d[319-260] ^ d[319-258] ^ d[319-256] ^ d[319-250] ^ d[319-249] ^ d[319-247] ^ d[319-244] ^ d[319-243] ^ d[319-240] ^ d[319-239] ^ d[319-236] ^ d[319-235] ^ d[319-229] ^ d[319-226] ^ d[319-225] ^ d[319-224] ^ d[319-223] ^ d[319-222] ^ d[319-220] ^ d[319-218] ^ d[319-217] ^ d[319-216] ^ d[319-211] ^ d[319-210] ^ d[319-209] ^ d[319-208] ^ d[319-204] ^ d[319-198] ^ d[319-197] ^ d[319-194] ^ d[319-193] ^ d[319-192] ^ d[319-191] ^ d[319-190] ^ d[319-187] ^ d[319-184] ^ d[319-183] ^ d[319-180] ^ d[319-179] ^ d[319-178] ^ d[319-175] ^ d[319-173] ^ d[319-171] ^ d[319-168] ^ d[319-165] ^ d[319-164] ^ d[319-163] ^ d[319-161] ^ d[319-160] ^ d[319-159] ^ d[319-157] ^ d[319-154] ^ d[319-153] ^ d[319-152] ^ d[319-151] ^ d[319-150] ^ d[319-149] ^ d[319-148] ^ d[319-141] ^ d[319-139] ^ d[319-136] ^ d[319-135] ^ d[319-134] ^ d[319-130] ^ d[319-127] ^ d[319-126] ^ d[319-125] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-117] ^ d[319-115] ^ d[319-113] ^ d[319-110] ^ d[319-109] ^ d[319-107] ^ d[319-106] ^ d[319-105] ^ d[319-104] ^ d[319-101] ^ d[319-98] ^ d[319-96] ^ d[319-95] ^ d[319-94] ^ d[319-90] ^ d[319-89] ^ d[319-86] ^ d[319-83] ^ d[319-80] ^ d[319-78] ^ d[319-77] ^ d[319-75] ^ d[319-73] ^ d[319-71] ^ d[319-70] ^ d[319-69] ^ d[319-66] ^ d[319-63] ^ d[319-62] ^ d[319-60] ^ d[319-59] ^ d[319-58] ^ d[319-56] ^ d[319-55] ^ d[319-52] ^ d[319-50] ^ d[319-42] ^ d[319-40] ^ d[319-39] ^ d[319-36] ^ d[319-35] ^ d[319-33] ^ d[319-32] ^ d[319-31] ^ d[319-29] ^ d[319-28] ^ d[319-26] ^ d[319-19] ^ d[319-16] ^ d[319-14] ^ d[319-13] ^ d[319-9] ^ d[319-5] ^ d[319-3] ^ d[319-2] ^ d[319-0] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-7] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-18] ^ c[31-19] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-30];
                stage_crc320_crc[20] <= d[319-318] ^ d[319-316] ^ d[319-314] ^ d[319-313] ^ d[319-312] ^ d[319-310] ^ d[319-309] ^ d[319-308] ^ d[319-307] ^ d[319-305] ^ d[319-301] ^ d[319-299] ^ d[319-298] ^ d[319-297] ^ d[319-295] ^ d[319-294] ^ d[319-293] ^ d[319-291] ^ d[319-290] ^ d[319-287] ^ d[319-286] ^ d[319-285] ^ d[319-282] ^ d[319-279] ^ d[319-277] ^ d[319-275] ^ d[319-274] ^ d[319-273] ^ d[319-267] ^ d[319-265] ^ d[319-263] ^ d[319-255] ^ d[319-252] ^ d[319-251] ^ d[319-250] ^ d[319-245] ^ d[319-244] ^ d[319-243] ^ d[319-241] ^ d[319-240] ^ d[319-236] ^ d[319-234] ^ d[319-228] ^ d[319-225] ^ d[319-223] ^ d[319-221] ^ d[319-219] ^ d[319-218] ^ d[319-217] ^ d[319-216] ^ d[319-214] ^ d[319-211] ^ d[319-208] ^ d[319-207] ^ d[319-205] ^ d[319-203] ^ d[319-202] ^ d[319-201] ^ d[319-197] ^ d[319-195] ^ d[319-190] ^ d[319-186] ^ d[319-185] ^ d[319-184] ^ d[319-183] ^ d[319-182] ^ d[319-181] ^ d[319-180] ^ d[319-179] ^ d[319-176] ^ d[319-174] ^ d[319-171] ^ d[319-170] ^ d[319-167] ^ d[319-165] ^ d[319-164] ^ d[319-160] ^ d[319-156] ^ d[319-154] ^ d[319-153] ^ d[319-152] ^ d[319-150] ^ d[319-144] ^ d[319-143] ^ d[319-142] ^ d[319-140] ^ d[319-134] ^ d[319-132] ^ d[319-131] ^ d[319-125] ^ d[319-124] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-117] ^ d[319-113] ^ d[319-108] ^ d[319-107] ^ d[319-105] ^ d[319-104] ^ d[319-103] ^ d[319-102] ^ d[319-101] ^ d[319-98] ^ d[319-94] ^ d[319-91] ^ d[319-90] ^ d[319-85] ^ d[319-83] ^ d[319-82] ^ d[319-78] ^ d[319-76] ^ d[319-74] ^ d[319-73] ^ d[319-71] ^ d[319-70] ^ d[319-68] ^ d[319-66] ^ d[319-65] ^ d[319-64] ^ d[319-59] ^ d[319-58] ^ d[319-57] ^ d[319-56] ^ d[319-55] ^ d[319-54] ^ d[319-51] ^ d[319-50] ^ d[319-48] ^ d[319-47] ^ d[319-45] ^ d[319-44] ^ d[319-43] ^ d[319-41] ^ d[319-40] ^ d[319-36] ^ d[319-33] ^ d[319-31] ^ d[319-28] ^ d[319-27] ^ d[319-26] ^ d[319-25] ^ d[319-24] ^ d[319-20] ^ d[319-17] ^ d[319-16] ^ d[319-15] ^ d[319-14] ^ d[319-12] ^ d[319-9] ^ d[319-4] ^ d[319-3] ^ d[319-1] ^ d[319-0] ^ c[31-2] ^ c[31-3] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-13] ^ c[31-17] ^ c[31-19] ^ c[31-20] ^ c[31-21] ^ c[31-22] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-28] ^ c[31-30];
                stage_crc320_crc[19] <= d[319-318] ^ d[319-314] ^ d[319-313] ^ d[319-312] ^ d[319-311] ^ d[319-308] ^ d[319-306] ^ d[319-305] ^ d[319-303] ^ d[319-297] ^ d[319-291] ^ d[319-290] ^ d[319-280] ^ d[319-279] ^ d[319-278] ^ d[319-277] ^ d[319-275] ^ d[319-273] ^ d[319-269] ^ d[319-266] ^ d[319-265] ^ d[319-261] ^ d[319-259] ^ d[319-257] ^ d[319-256] ^ d[319-255] ^ d[319-253] ^ d[319-251] ^ d[319-248] ^ d[319-246] ^ d[319-245] ^ d[319-244] ^ d[319-243] ^ d[319-242] ^ d[319-241] ^ d[319-235] ^ d[319-234] ^ d[319-230] ^ d[319-229] ^ d[319-228] ^ d[319-227] ^ d[319-222] ^ d[319-220] ^ d[319-219] ^ d[319-218] ^ d[319-217] ^ d[319-216] ^ d[319-215] ^ d[319-214] ^ d[319-210] ^ d[319-207] ^ d[319-206] ^ d[319-204] ^ d[319-201] ^ d[319-199] ^ d[319-197] ^ d[319-196] ^ d[319-194] ^ d[319-193] ^ d[319-192] ^ d[319-190] ^ d[319-188] ^ d[319-187] ^ d[319-185] ^ d[319-184] ^ d[319-181] ^ d[319-180] ^ d[319-177] ^ d[319-175] ^ d[319-170] ^ d[319-169] ^ d[319-168] ^ d[319-167] ^ d[319-165] ^ d[319-162] ^ d[319-158] ^ d[319-157] ^ d[319-156] ^ d[319-154] ^ d[319-153] ^ d[319-149] ^ d[319-145] ^ d[319-141] ^ d[319-137] ^ d[319-136] ^ d[319-134] ^ d[319-133] ^ d[319-128] ^ d[319-127] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-117] ^ d[319-116] ^ d[319-113] ^ d[319-111] ^ d[319-110] ^ d[319-109] ^ d[319-108] ^ d[319-105] ^ d[319-102] ^ d[319-101] ^ d[319-98] ^ d[319-97] ^ d[319-96] ^ d[319-94] ^ d[319-92] ^ d[319-91] ^ d[319-87] ^ d[319-86] ^ d[319-85] ^ d[319-82] ^ d[319-81] ^ d[319-77] ^ d[319-75] ^ d[319-74] ^ d[319-73] ^ d[319-71] ^ d[319-69] ^ d[319-68] ^ d[319-63] ^ d[319-61] ^ d[319-59] ^ d[319-57] ^ d[319-56] ^ d[319-54] ^ d[319-53] ^ d[319-52] ^ d[319-51] ^ d[319-50] ^ d[319-49] ^ d[319-47] ^ d[319-46] ^ d[319-42] ^ d[319-41] ^ d[319-31] ^ d[319-30] ^ d[319-27] ^ d[319-24] ^ d[319-21] ^ d[319-18] ^ d[319-17] ^ d[319-15] ^ d[319-13] ^ d[319-12] ^ d[319-9] ^ d[319-6] ^ d[319-5] ^ d[319-4] ^ d[319-2] ^ d[319-1] ^ d[319-0] ^ c[31-2] ^ c[31-3] ^ c[31-9] ^ c[31-15] ^ c[31-17] ^ c[31-18] ^ c[31-20] ^ c[31-23] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-30];
                stage_crc320_crc[18] <= d[319-319] ^ d[319-315] ^ d[319-314] ^ d[319-313] ^ d[319-312] ^ d[319-309] ^ d[319-307] ^ d[319-306] ^ d[319-304] ^ d[319-298] ^ d[319-292] ^ d[319-291] ^ d[319-281] ^ d[319-280] ^ d[319-279] ^ d[319-278] ^ d[319-276] ^ d[319-274] ^ d[319-270] ^ d[319-267] ^ d[319-266] ^ d[319-262] ^ d[319-260] ^ d[319-258] ^ d[319-257] ^ d[319-256] ^ d[319-254] ^ d[319-252] ^ d[319-249] ^ d[319-247] ^ d[319-246] ^ d[319-245] ^ d[319-244] ^ d[319-243] ^ d[319-242] ^ d[319-236] ^ d[319-235] ^ d[319-231] ^ d[319-230] ^ d[319-229] ^ d[319-228] ^ d[319-223] ^ d[319-221] ^ d[319-220] ^ d[319-219] ^ d[319-218] ^ d[319-217] ^ d[319-216] ^ d[319-215] ^ d[319-211] ^ d[319-208] ^ d[319-207] ^ d[319-205] ^ d[319-202] ^ d[319-200] ^ d[319-198] ^ d[319-197] ^ d[319-195] ^ d[319-194] ^ d[319-193] ^ d[319-191] ^ d[319-189] ^ d[319-188] ^ d[319-186] ^ d[319-185] ^ d[319-182] ^ d[319-181] ^ d[319-178] ^ d[319-176] ^ d[319-171] ^ d[319-170] ^ d[319-169] ^ d[319-168] ^ d[319-166] ^ d[319-163] ^ d[319-159] ^ d[319-158] ^ d[319-157] ^ d[319-155] ^ d[319-154] ^ d[319-150] ^ d[319-146] ^ d[319-142] ^ d[319-138] ^ d[319-137] ^ d[319-135] ^ d[319-134] ^ d[319-129] ^ d[319-128] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-118] ^ d[319-117] ^ d[319-114] ^ d[319-112] ^ d[319-111] ^ d[319-110] ^ d[319-109] ^ d[319-106] ^ d[319-103] ^ d[319-102] ^ d[319-99] ^ d[319-98] ^ d[319-97] ^ d[319-95] ^ d[319-93] ^ d[319-92] ^ d[319-88] ^ d[319-87] ^ d[319-86] ^ d[319-83] ^ d[319-82] ^ d[319-78] ^ d[319-76] ^ d[319-75] ^ d[319-74] ^ d[319-72] ^ d[319-70] ^ d[319-69] ^ d[319-64] ^ d[319-62] ^ d[319-60] ^ d[319-58] ^ d[319-57] ^ d[319-55] ^ d[319-54] ^ d[319-53] ^ d[319-52] ^ d[319-51] ^ d[319-50] ^ d[319-48] ^ d[319-47] ^ d[319-43] ^ d[319-42] ^ d[319-32] ^ d[319-31] ^ d[319-28] ^ d[319-25] ^ d[319-22] ^ d[319-19] ^ d[319-18] ^ d[319-16] ^ d[319-14] ^ d[319-13] ^ d[319-10] ^ d[319-7] ^ d[319-6] ^ d[319-5] ^ d[319-3] ^ d[319-2] ^ d[319-1] ^ c[31-3] ^ c[31-4] ^ c[31-10] ^ c[31-16] ^ c[31-18] ^ c[31-19] ^ c[31-21] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-31];
                stage_crc320_crc[17] <= d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-313] ^ d[319-310] ^ d[319-308] ^ d[319-307] ^ d[319-305] ^ d[319-299] ^ d[319-293] ^ d[319-292] ^ d[319-282] ^ d[319-281] ^ d[319-280] ^ d[319-279] ^ d[319-277] ^ d[319-275] ^ d[319-271] ^ d[319-268] ^ d[319-267] ^ d[319-263] ^ d[319-261] ^ d[319-259] ^ d[319-258] ^ d[319-257] ^ d[319-255] ^ d[319-253] ^ d[319-250] ^ d[319-248] ^ d[319-247] ^ d[319-246] ^ d[319-245] ^ d[319-244] ^ d[319-243] ^ d[319-237] ^ d[319-236] ^ d[319-232] ^ d[319-231] ^ d[319-230] ^ d[319-229] ^ d[319-224] ^ d[319-222] ^ d[319-221] ^ d[319-220] ^ d[319-219] ^ d[319-218] ^ d[319-217] ^ d[319-216] ^ d[319-212] ^ d[319-209] ^ d[319-208] ^ d[319-206] ^ d[319-203] ^ d[319-201] ^ d[319-199] ^ d[319-198] ^ d[319-196] ^ d[319-195] ^ d[319-194] ^ d[319-192] ^ d[319-190] ^ d[319-189] ^ d[319-187] ^ d[319-186] ^ d[319-183] ^ d[319-182] ^ d[319-179] ^ d[319-177] ^ d[319-172] ^ d[319-171] ^ d[319-170] ^ d[319-169] ^ d[319-167] ^ d[319-164] ^ d[319-160] ^ d[319-159] ^ d[319-158] ^ d[319-156] ^ d[319-155] ^ d[319-151] ^ d[319-147] ^ d[319-143] ^ d[319-139] ^ d[319-138] ^ d[319-136] ^ d[319-135] ^ d[319-130] ^ d[319-129] ^ d[319-124] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-119] ^ d[319-118] ^ d[319-115] ^ d[319-113] ^ d[319-112] ^ d[319-111] ^ d[319-110] ^ d[319-107] ^ d[319-104] ^ d[319-103] ^ d[319-100] ^ d[319-99] ^ d[319-98] ^ d[319-96] ^ d[319-94] ^ d[319-93] ^ d[319-89] ^ d[319-88] ^ d[319-87] ^ d[319-84] ^ d[319-83] ^ d[319-79] ^ d[319-77] ^ d[319-76] ^ d[319-75] ^ d[319-73] ^ d[319-71] ^ d[319-70] ^ d[319-65] ^ d[319-63] ^ d[319-61] ^ d[319-59] ^ d[319-58] ^ d[319-56] ^ d[319-55] ^ d[319-54] ^ d[319-53] ^ d[319-52] ^ d[319-51] ^ d[319-49] ^ d[319-48] ^ d[319-44] ^ d[319-43] ^ d[319-33] ^ d[319-32] ^ d[319-29] ^ d[319-26] ^ d[319-23] ^ d[319-20] ^ d[319-19] ^ d[319-17] ^ d[319-15] ^ d[319-14] ^ d[319-11] ^ d[319-8] ^ d[319-7] ^ d[319-6] ^ d[319-4] ^ d[319-3] ^ d[319-2] ^ c[31-4] ^ c[31-5] ^ c[31-11] ^ c[31-17] ^ c[31-19] ^ c[31-20] ^ c[31-22] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28];
                stage_crc320_crc[16] <= d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-311] ^ d[319-309] ^ d[319-308] ^ d[319-306] ^ d[319-300] ^ d[319-294] ^ d[319-293] ^ d[319-283] ^ d[319-282] ^ d[319-281] ^ d[319-280] ^ d[319-278] ^ d[319-276] ^ d[319-272] ^ d[319-269] ^ d[319-268] ^ d[319-264] ^ d[319-262] ^ d[319-260] ^ d[319-259] ^ d[319-258] ^ d[319-256] ^ d[319-254] ^ d[319-251] ^ d[319-249] ^ d[319-248] ^ d[319-247] ^ d[319-246] ^ d[319-245] ^ d[319-244] ^ d[319-238] ^ d[319-237] ^ d[319-233] ^ d[319-232] ^ d[319-231] ^ d[319-230] ^ d[319-225] ^ d[319-223] ^ d[319-222] ^ d[319-221] ^ d[319-220] ^ d[319-219] ^ d[319-218] ^ d[319-217] ^ d[319-213] ^ d[319-210] ^ d[319-209] ^ d[319-207] ^ d[319-204] ^ d[319-202] ^ d[319-200] ^ d[319-199] ^ d[319-197] ^ d[319-196] ^ d[319-195] ^ d[319-193] ^ d[319-191] ^ d[319-190] ^ d[319-188] ^ d[319-187] ^ d[319-184] ^ d[319-183] ^ d[319-180] ^ d[319-178] ^ d[319-173] ^ d[319-172] ^ d[319-171] ^ d[319-170] ^ d[319-168] ^ d[319-165] ^ d[319-161] ^ d[319-160] ^ d[319-159] ^ d[319-157] ^ d[319-156] ^ d[319-152] ^ d[319-148] ^ d[319-144] ^ d[319-140] ^ d[319-139] ^ d[319-137] ^ d[319-136] ^ d[319-131] ^ d[319-130] ^ d[319-125] ^ d[319-124] ^ d[319-123] ^ d[319-122] ^ d[319-120] ^ d[319-119] ^ d[319-116] ^ d[319-114] ^ d[319-113] ^ d[319-112] ^ d[319-111] ^ d[319-108] ^ d[319-105] ^ d[319-104] ^ d[319-101] ^ d[319-100] ^ d[319-99] ^ d[319-97] ^ d[319-95] ^ d[319-94] ^ d[319-90] ^ d[319-89] ^ d[319-88] ^ d[319-85] ^ d[319-84] ^ d[319-80] ^ d[319-78] ^ d[319-77] ^ d[319-76] ^ d[319-74] ^ d[319-72] ^ d[319-71] ^ d[319-66] ^ d[319-64] ^ d[319-62] ^ d[319-60] ^ d[319-59] ^ d[319-57] ^ d[319-56] ^ d[319-55] ^ d[319-54] ^ d[319-53] ^ d[319-52] ^ d[319-50] ^ d[319-49] ^ d[319-45] ^ d[319-44] ^ d[319-34] ^ d[319-33] ^ d[319-30] ^ d[319-27] ^ d[319-24] ^ d[319-21] ^ d[319-20] ^ d[319-18] ^ d[319-16] ^ d[319-15] ^ d[319-12] ^ d[319-9] ^ d[319-8] ^ d[319-7] ^ d[319-5] ^ d[319-4] ^ d[319-3] ^ c[31-5] ^ c[31-6] ^ c[31-12] ^ c[31-18] ^ c[31-20] ^ c[31-21] ^ c[31-23] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29];
                stage_crc320_crc[15] <= d[319-319] ^ d[319-316] ^ d[319-307] ^ d[319-305] ^ d[319-303] ^ d[319-302] ^ d[319-301] ^ d[319-300] ^ d[319-299] ^ d[319-298] ^ d[319-297] ^ d[319-296] ^ d[319-292] ^ d[319-290] ^ d[319-288] ^ d[319-287] ^ d[319-286] ^ d[319-284] ^ d[319-282] ^ d[319-281] ^ d[319-276] ^ d[319-274] ^ d[319-270] ^ d[319-268] ^ d[319-264] ^ d[319-263] ^ d[319-260] ^ d[319-250] ^ d[319-249] ^ d[319-247] ^ d[319-246] ^ d[319-245] ^ d[319-243] ^ d[319-239] ^ d[319-238] ^ d[319-237] ^ d[319-233] ^ d[319-232] ^ d[319-231] ^ d[319-230] ^ d[319-228] ^ d[319-227] ^ d[319-223] ^ d[319-222] ^ d[319-221] ^ d[319-220] ^ d[319-219] ^ d[319-218] ^ d[319-216] ^ d[319-212] ^ d[319-211] ^ d[319-209] ^ d[319-207] ^ d[319-205] ^ d[319-202] ^ d[319-200] ^ d[319-199] ^ d[319-196] ^ d[319-193] ^ d[319-190] ^ d[319-189] ^ d[319-186] ^ d[319-185] ^ d[319-184] ^ d[319-183] ^ d[319-182] ^ d[319-181] ^ d[319-179] ^ d[319-174] ^ d[319-173] ^ d[319-170] ^ d[319-167] ^ d[319-160] ^ d[319-157] ^ d[319-156] ^ d[319-155] ^ d[319-153] ^ d[319-151] ^ d[319-145] ^ d[319-144] ^ d[319-143] ^ d[319-141] ^ d[319-140] ^ d[319-138] ^ d[319-136] ^ d[319-135] ^ d[319-134] ^ d[319-131] ^ d[319-128] ^ d[319-127] ^ d[319-124] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-118] ^ d[319-116] ^ d[319-115] ^ d[319-112] ^ d[319-111] ^ d[319-110] ^ d[319-109] ^ d[319-105] ^ d[319-104] ^ d[319-103] ^ d[319-102] ^ d[319-100] ^ d[319-99] ^ d[319-97] ^ d[319-94] ^ d[319-91] ^ d[319-90] ^ d[319-89] ^ d[319-87] ^ d[319-86] ^ d[319-84] ^ d[319-83] ^ d[319-82] ^ d[319-78] ^ d[319-77] ^ d[319-75] ^ d[319-68] ^ d[319-66] ^ d[319-57] ^ d[319-56] ^ d[319-51] ^ d[319-48] ^ d[319-47] ^ d[319-46] ^ d[319-44] ^ d[319-37] ^ d[319-35] ^ d[319-32] ^ d[319-30] ^ d[319-29] ^ d[319-26] ^ d[319-24] ^ d[319-22] ^ d[319-21] ^ d[319-19] ^ d[319-17] ^ d[319-13] ^ d[319-12] ^ d[319-8] ^ d[319-5] ^ d[319-4] ^ d[319-0] ^ c[31-0] ^ c[31-2] ^ c[31-4] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-17] ^ c[31-19] ^ c[31-28] ^ c[31-31];
                stage_crc320_crc[14] <= d[319-317] ^ d[319-308] ^ d[319-306] ^ d[319-304] ^ d[319-303] ^ d[319-302] ^ d[319-301] ^ d[319-300] ^ d[319-299] ^ d[319-298] ^ d[319-297] ^ d[319-293] ^ d[319-291] ^ d[319-289] ^ d[319-288] ^ d[319-287] ^ d[319-285] ^ d[319-283] ^ d[319-282] ^ d[319-277] ^ d[319-275] ^ d[319-271] ^ d[319-269] ^ d[319-265] ^ d[319-264] ^ d[319-261] ^ d[319-251] ^ d[319-250] ^ d[319-248] ^ d[319-247] ^ d[319-246] ^ d[319-244] ^ d[319-240] ^ d[319-239] ^ d[319-238] ^ d[319-234] ^ d[319-233] ^ d[319-232] ^ d[319-231] ^ d[319-229] ^ d[319-228] ^ d[319-224] ^ d[319-223] ^ d[319-222] ^ d[319-221] ^ d[319-220] ^ d[319-219] ^ d[319-217] ^ d[319-213] ^ d[319-212] ^ d[319-210] ^ d[319-208] ^ d[319-206] ^ d[319-203] ^ d[319-201] ^ d[319-200] ^ d[319-197] ^ d[319-194] ^ d[319-191] ^ d[319-190] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-184] ^ d[319-183] ^ d[319-182] ^ d[319-180] ^ d[319-175] ^ d[319-174] ^ d[319-171] ^ d[319-168] ^ d[319-161] ^ d[319-158] ^ d[319-157] ^ d[319-156] ^ d[319-154] ^ d[319-152] ^ d[319-146] ^ d[319-145] ^ d[319-144] ^ d[319-142] ^ d[319-141] ^ d[319-139] ^ d[319-137] ^ d[319-136] ^ d[319-135] ^ d[319-132] ^ d[319-129] ^ d[319-128] ^ d[319-125] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-117] ^ d[319-116] ^ d[319-113] ^ d[319-112] ^ d[319-111] ^ d[319-110] ^ d[319-106] ^ d[319-105] ^ d[319-104] ^ d[319-103] ^ d[319-101] ^ d[319-100] ^ d[319-98] ^ d[319-95] ^ d[319-92] ^ d[319-91] ^ d[319-90] ^ d[319-88] ^ d[319-87] ^ d[319-85] ^ d[319-84] ^ d[319-83] ^ d[319-79] ^ d[319-78] ^ d[319-76] ^ d[319-69] ^ d[319-67] ^ d[319-58] ^ d[319-57] ^ d[319-52] ^ d[319-49] ^ d[319-48] ^ d[319-47] ^ d[319-45] ^ d[319-38] ^ d[319-36] ^ d[319-33] ^ d[319-31] ^ d[319-30] ^ d[319-27] ^ d[319-25] ^ d[319-23] ^ d[319-22] ^ d[319-20] ^ d[319-18] ^ d[319-14] ^ d[319-13] ^ d[319-9] ^ d[319-6] ^ d[319-5] ^ d[319-1] ^ c[31-0] ^ c[31-1] ^ c[31-3] ^ c[31-5] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-18] ^ c[31-20] ^ c[31-29];
                stage_crc320_crc[13] <= d[319-318] ^ d[319-309] ^ d[319-307] ^ d[319-305] ^ d[319-304] ^ d[319-303] ^ d[319-302] ^ d[319-301] ^ d[319-300] ^ d[319-299] ^ d[319-298] ^ d[319-294] ^ d[319-292] ^ d[319-290] ^ d[319-289] ^ d[319-288] ^ d[319-286] ^ d[319-284] ^ d[319-283] ^ d[319-278] ^ d[319-276] ^ d[319-272] ^ d[319-270] ^ d[319-266] ^ d[319-265] ^ d[319-262] ^ d[319-252] ^ d[319-251] ^ d[319-249] ^ d[319-248] ^ d[319-247] ^ d[319-245] ^ d[319-241] ^ d[319-240] ^ d[319-239] ^ d[319-235] ^ d[319-234] ^ d[319-233] ^ d[319-232] ^ d[319-230] ^ d[319-229] ^ d[319-225] ^ d[319-224] ^ d[319-223] ^ d[319-222] ^ d[319-221] ^ d[319-220] ^ d[319-218] ^ d[319-214] ^ d[319-213] ^ d[319-211] ^ d[319-209] ^ d[319-207] ^ d[319-204] ^ d[319-202] ^ d[319-201] ^ d[319-198] ^ d[319-195] ^ d[319-192] ^ d[319-191] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-184] ^ d[319-183] ^ d[319-181] ^ d[319-176] ^ d[319-175] ^ d[319-172] ^ d[319-169] ^ d[319-162] ^ d[319-159] ^ d[319-158] ^ d[319-157] ^ d[319-155] ^ d[319-153] ^ d[319-147] ^ d[319-146] ^ d[319-145] ^ d[319-143] ^ d[319-142] ^ d[319-140] ^ d[319-138] ^ d[319-137] ^ d[319-136] ^ d[319-133] ^ d[319-130] ^ d[319-129] ^ d[319-126] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-118] ^ d[319-117] ^ d[319-114] ^ d[319-113] ^ d[319-112] ^ d[319-111] ^ d[319-107] ^ d[319-106] ^ d[319-105] ^ d[319-104] ^ d[319-102] ^ d[319-101] ^ d[319-99] ^ d[319-96] ^ d[319-93] ^ d[319-92] ^ d[319-91] ^ d[319-89] ^ d[319-88] ^ d[319-86] ^ d[319-85] ^ d[319-84] ^ d[319-80] ^ d[319-79] ^ d[319-77] ^ d[319-70] ^ d[319-68] ^ d[319-59] ^ d[319-58] ^ d[319-53] ^ d[319-50] ^ d[319-49] ^ d[319-48] ^ d[319-46] ^ d[319-39] ^ d[319-37] ^ d[319-34] ^ d[319-32] ^ d[319-31] ^ d[319-28] ^ d[319-26] ^ d[319-24] ^ d[319-23] ^ d[319-21] ^ d[319-19] ^ d[319-15] ^ d[319-14] ^ d[319-10] ^ d[319-7] ^ d[319-6] ^ d[319-2] ^ c[31-0] ^ c[31-1] ^ c[31-2] ^ c[31-4] ^ c[31-6] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-19] ^ c[31-21] ^ c[31-30];
                stage_crc320_crc[12] <= d[319-319] ^ d[319-310] ^ d[319-308] ^ d[319-306] ^ d[319-305] ^ d[319-304] ^ d[319-303] ^ d[319-302] ^ d[319-301] ^ d[319-300] ^ d[319-299] ^ d[319-295] ^ d[319-293] ^ d[319-291] ^ d[319-290] ^ d[319-289] ^ d[319-287] ^ d[319-285] ^ d[319-284] ^ d[319-279] ^ d[319-277] ^ d[319-273] ^ d[319-271] ^ d[319-267] ^ d[319-266] ^ d[319-263] ^ d[319-253] ^ d[319-252] ^ d[319-250] ^ d[319-249] ^ d[319-248] ^ d[319-246] ^ d[319-242] ^ d[319-241] ^ d[319-240] ^ d[319-236] ^ d[319-235] ^ d[319-234] ^ d[319-233] ^ d[319-231] ^ d[319-230] ^ d[319-226] ^ d[319-225] ^ d[319-224] ^ d[319-223] ^ d[319-222] ^ d[319-221] ^ d[319-219] ^ d[319-215] ^ d[319-214] ^ d[319-212] ^ d[319-210] ^ d[319-208] ^ d[319-205] ^ d[319-203] ^ d[319-202] ^ d[319-199] ^ d[319-196] ^ d[319-193] ^ d[319-192] ^ d[319-189] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-184] ^ d[319-182] ^ d[319-177] ^ d[319-176] ^ d[319-173] ^ d[319-170] ^ d[319-163] ^ d[319-160] ^ d[319-159] ^ d[319-158] ^ d[319-156] ^ d[319-154] ^ d[319-148] ^ d[319-147] ^ d[319-146] ^ d[319-144] ^ d[319-143] ^ d[319-141] ^ d[319-139] ^ d[319-138] ^ d[319-137] ^ d[319-134] ^ d[319-131] ^ d[319-130] ^ d[319-127] ^ d[319-124] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-119] ^ d[319-118] ^ d[319-115] ^ d[319-114] ^ d[319-113] ^ d[319-112] ^ d[319-108] ^ d[319-107] ^ d[319-106] ^ d[319-105] ^ d[319-103] ^ d[319-102] ^ d[319-100] ^ d[319-97] ^ d[319-94] ^ d[319-93] ^ d[319-92] ^ d[319-90] ^ d[319-89] ^ d[319-87] ^ d[319-86] ^ d[319-85] ^ d[319-81] ^ d[319-80] ^ d[319-78] ^ d[319-71] ^ d[319-69] ^ d[319-60] ^ d[319-59] ^ d[319-54] ^ d[319-51] ^ d[319-50] ^ d[319-49] ^ d[319-47] ^ d[319-40] ^ d[319-38] ^ d[319-35] ^ d[319-33] ^ d[319-32] ^ d[319-29] ^ d[319-27] ^ d[319-25] ^ d[319-24] ^ d[319-22] ^ d[319-20] ^ d[319-16] ^ d[319-15] ^ d[319-11] ^ d[319-8] ^ d[319-7] ^ d[319-3] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-5] ^ c[31-7] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-20] ^ c[31-22] ^ c[31-31];
                stage_crc320_crc[11] <= d[319-311] ^ d[319-309] ^ d[319-307] ^ d[319-306] ^ d[319-305] ^ d[319-304] ^ d[319-303] ^ d[319-302] ^ d[319-301] ^ d[319-300] ^ d[319-296] ^ d[319-294] ^ d[319-292] ^ d[319-291] ^ d[319-290] ^ d[319-288] ^ d[319-286] ^ d[319-285] ^ d[319-280] ^ d[319-278] ^ d[319-274] ^ d[319-272] ^ d[319-268] ^ d[319-267] ^ d[319-264] ^ d[319-254] ^ d[319-253] ^ d[319-251] ^ d[319-250] ^ d[319-249] ^ d[319-247] ^ d[319-243] ^ d[319-242] ^ d[319-241] ^ d[319-237] ^ d[319-236] ^ d[319-235] ^ d[319-234] ^ d[319-232] ^ d[319-231] ^ d[319-227] ^ d[319-226] ^ d[319-225] ^ d[319-224] ^ d[319-223] ^ d[319-222] ^ d[319-220] ^ d[319-216] ^ d[319-215] ^ d[319-213] ^ d[319-211] ^ d[319-209] ^ d[319-206] ^ d[319-204] ^ d[319-203] ^ d[319-200] ^ d[319-197] ^ d[319-194] ^ d[319-193] ^ d[319-190] ^ d[319-189] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-183] ^ d[319-178] ^ d[319-177] ^ d[319-174] ^ d[319-171] ^ d[319-164] ^ d[319-161] ^ d[319-160] ^ d[319-159] ^ d[319-157] ^ d[319-155] ^ d[319-149] ^ d[319-148] ^ d[319-147] ^ d[319-145] ^ d[319-144] ^ d[319-142] ^ d[319-140] ^ d[319-139] ^ d[319-138] ^ d[319-135] ^ d[319-132] ^ d[319-131] ^ d[319-128] ^ d[319-125] ^ d[319-124] ^ d[319-123] ^ d[319-122] ^ d[319-120] ^ d[319-119] ^ d[319-116] ^ d[319-115] ^ d[319-114] ^ d[319-113] ^ d[319-109] ^ d[319-108] ^ d[319-107] ^ d[319-106] ^ d[319-104] ^ d[319-103] ^ d[319-101] ^ d[319-98] ^ d[319-95] ^ d[319-94] ^ d[319-93] ^ d[319-91] ^ d[319-90] ^ d[319-88] ^ d[319-87] ^ d[319-86] ^ d[319-82] ^ d[319-81] ^ d[319-79] ^ d[319-72] ^ d[319-70] ^ d[319-61] ^ d[319-60] ^ d[319-55] ^ d[319-52] ^ d[319-51] ^ d[319-50] ^ d[319-48] ^ d[319-41] ^ d[319-39] ^ d[319-36] ^ d[319-34] ^ d[319-33] ^ d[319-30] ^ d[319-28] ^ d[319-26] ^ d[319-25] ^ d[319-23] ^ d[319-21] ^ d[319-17] ^ d[319-16] ^ d[319-12] ^ d[319-9] ^ d[319-8] ^ d[319-4] ^ c[31-0] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-6] ^ c[31-8] ^ c[31-12] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-19] ^ c[31-21] ^ c[31-23];
                stage_crc320_crc[10] <= d[319-312] ^ d[319-310] ^ d[319-308] ^ d[319-307] ^ d[319-306] ^ d[319-305] ^ d[319-304] ^ d[319-303] ^ d[319-302] ^ d[319-301] ^ d[319-297] ^ d[319-295] ^ d[319-293] ^ d[319-292] ^ d[319-291] ^ d[319-289] ^ d[319-287] ^ d[319-286] ^ d[319-281] ^ d[319-279] ^ d[319-275] ^ d[319-273] ^ d[319-269] ^ d[319-268] ^ d[319-265] ^ d[319-255] ^ d[319-254] ^ d[319-252] ^ d[319-251] ^ d[319-250] ^ d[319-248] ^ d[319-244] ^ d[319-243] ^ d[319-242] ^ d[319-238] ^ d[319-237] ^ d[319-236] ^ d[319-235] ^ d[319-233] ^ d[319-232] ^ d[319-228] ^ d[319-227] ^ d[319-226] ^ d[319-225] ^ d[319-224] ^ d[319-223] ^ d[319-221] ^ d[319-217] ^ d[319-216] ^ d[319-214] ^ d[319-212] ^ d[319-210] ^ d[319-207] ^ d[319-205] ^ d[319-204] ^ d[319-201] ^ d[319-198] ^ d[319-195] ^ d[319-194] ^ d[319-191] ^ d[319-190] ^ d[319-189] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-184] ^ d[319-179] ^ d[319-178] ^ d[319-175] ^ d[319-172] ^ d[319-165] ^ d[319-162] ^ d[319-161] ^ d[319-160] ^ d[319-158] ^ d[319-156] ^ d[319-150] ^ d[319-149] ^ d[319-148] ^ d[319-146] ^ d[319-145] ^ d[319-143] ^ d[319-141] ^ d[319-140] ^ d[319-139] ^ d[319-136] ^ d[319-133] ^ d[319-132] ^ d[319-129] ^ d[319-126] ^ d[319-125] ^ d[319-124] ^ d[319-123] ^ d[319-121] ^ d[319-120] ^ d[319-117] ^ d[319-116] ^ d[319-115] ^ d[319-114] ^ d[319-110] ^ d[319-109] ^ d[319-108] ^ d[319-107] ^ d[319-105] ^ d[319-104] ^ d[319-102] ^ d[319-99] ^ d[319-96] ^ d[319-95] ^ d[319-94] ^ d[319-92] ^ d[319-91] ^ d[319-89] ^ d[319-88] ^ d[319-87] ^ d[319-83] ^ d[319-82] ^ d[319-80] ^ d[319-73] ^ d[319-71] ^ d[319-62] ^ d[319-61] ^ d[319-56] ^ d[319-53] ^ d[319-52] ^ d[319-51] ^ d[319-49] ^ d[319-42] ^ d[319-40] ^ d[319-37] ^ d[319-35] ^ d[319-34] ^ d[319-31] ^ d[319-29] ^ d[319-27] ^ d[319-26] ^ d[319-24] ^ d[319-22] ^ d[319-18] ^ d[319-17] ^ d[319-13] ^ d[319-10] ^ d[319-9] ^ d[319-5] ^ c[31-1] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-7] ^ c[31-9] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-19] ^ c[31-20] ^ c[31-22] ^ c[31-24];
                stage_crc320_crc[9] <= d[319-319] ^ d[319-318] ^ d[319-317] ^ d[319-315] ^ d[319-313] ^ d[319-312] ^ d[319-311] ^ d[319-310] ^ d[319-308] ^ d[319-307] ^ d[319-306] ^ d[319-304] ^ d[319-300] ^ d[319-299] ^ d[319-297] ^ d[319-295] ^ d[319-293] ^ d[319-286] ^ d[319-283] ^ d[319-282] ^ d[319-280] ^ d[319-279] ^ d[319-277] ^ d[319-273] ^ d[319-270] ^ d[319-268] ^ d[319-266] ^ d[319-265] ^ d[319-264] ^ d[319-261] ^ d[319-259] ^ d[319-257] ^ d[319-256] ^ d[319-253] ^ d[319-251] ^ d[319-249] ^ d[319-248] ^ d[319-245] ^ d[319-244] ^ d[319-239] ^ d[319-238] ^ d[319-236] ^ d[319-233] ^ d[319-230] ^ d[319-229] ^ d[319-225] ^ d[319-222] ^ d[319-218] ^ d[319-217] ^ d[319-216] ^ d[319-215] ^ d[319-214] ^ d[319-213] ^ d[319-212] ^ d[319-211] ^ d[319-210] ^ d[319-209] ^ d[319-207] ^ d[319-206] ^ d[319-205] ^ d[319-203] ^ d[319-201] ^ d[319-198] ^ d[319-197] ^ d[319-196] ^ d[319-195] ^ d[319-194] ^ d[319-193] ^ d[319-189] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-183] ^ d[319-182] ^ d[319-180] ^ d[319-179] ^ d[319-176] ^ d[319-173] ^ d[319-172] ^ d[319-171] ^ d[319-170] ^ d[319-169] ^ d[319-167] ^ d[319-163] ^ d[319-159] ^ d[319-158] ^ d[319-157] ^ d[319-156] ^ d[319-155] ^ d[319-150] ^ d[319-147] ^ d[319-146] ^ d[319-143] ^ d[319-142] ^ d[319-141] ^ d[319-140] ^ d[319-136] ^ d[319-135] ^ d[319-133] ^ d[319-132] ^ d[319-130] ^ d[319-128] ^ d[319-124] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-119] ^ d[319-115] ^ d[319-114] ^ d[319-113] ^ d[319-109] ^ d[319-108] ^ d[319-105] ^ d[319-104] ^ d[319-101] ^ d[319-100] ^ d[319-99] ^ d[319-98] ^ d[319-94] ^ d[319-93] ^ d[319-92] ^ d[319-90] ^ d[319-89] ^ d[319-88] ^ d[319-87] ^ d[319-85] ^ d[319-82] ^ d[319-79] ^ d[319-74] ^ d[319-73] ^ d[319-68] ^ d[319-67] ^ d[319-66] ^ d[319-65] ^ d[319-62] ^ d[319-61] ^ d[319-60] ^ d[319-58] ^ d[319-57] ^ d[319-55] ^ d[319-52] ^ d[319-48] ^ d[319-47] ^ d[319-45] ^ d[319-44] ^ d[319-43] ^ d[319-41] ^ d[319-38] ^ d[319-37] ^ d[319-36] ^ d[319-35] ^ d[319-34] ^ d[319-31] ^ d[319-29] ^ d[319-27] ^ d[319-26] ^ d[319-24] ^ d[319-23] ^ d[319-19] ^ d[319-18] ^ d[319-16] ^ d[319-14] ^ d[319-12] ^ d[319-11] ^ d[319-9] ^ d[319-0] ^ c[31-5] ^ c[31-7] ^ c[31-9] ^ c[31-11] ^ c[31-12] ^ c[31-16] ^ c[31-18] ^ c[31-19] ^ c[31-20] ^ c[31-22] ^ c[31-23] ^ c[31-24] ^ c[31-25] ^ c[31-27] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc320_crc[8] <= d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-313] ^ d[319-311] ^ d[319-310] ^ d[319-308] ^ d[319-307] ^ d[319-303] ^ d[319-302] ^ d[319-301] ^ d[319-299] ^ d[319-297] ^ d[319-295] ^ d[319-292] ^ d[319-290] ^ d[319-288] ^ d[319-286] ^ d[319-284] ^ d[319-281] ^ d[319-280] ^ d[319-279] ^ d[319-278] ^ d[319-277] ^ d[319-276] ^ d[319-273] ^ d[319-271] ^ d[319-268] ^ d[319-267] ^ d[319-266] ^ d[319-264] ^ d[319-262] ^ d[319-261] ^ d[319-260] ^ d[319-259] ^ d[319-258] ^ d[319-255] ^ d[319-254] ^ d[319-250] ^ d[319-249] ^ d[319-248] ^ d[319-246] ^ d[319-245] ^ d[319-243] ^ d[319-240] ^ d[319-239] ^ d[319-231] ^ d[319-228] ^ d[319-227] ^ d[319-224] ^ d[319-223] ^ d[319-219] ^ d[319-218] ^ d[319-217] ^ d[319-215] ^ d[319-213] ^ d[319-211] ^ d[319-209] ^ d[319-206] ^ d[319-204] ^ d[319-203] ^ d[319-201] ^ d[319-196] ^ d[319-195] ^ d[319-193] ^ d[319-192] ^ d[319-191] ^ d[319-187] ^ d[319-184] ^ d[319-182] ^ d[319-181] ^ d[319-180] ^ d[319-177] ^ d[319-174] ^ d[319-173] ^ d[319-169] ^ d[319-168] ^ d[319-167] ^ d[319-166] ^ d[319-164] ^ d[319-162] ^ d[319-161] ^ d[319-160] ^ d[319-159] ^ d[319-157] ^ d[319-155] ^ d[319-149] ^ d[319-148] ^ d[319-147] ^ d[319-142] ^ d[319-141] ^ d[319-135] ^ d[319-133] ^ d[319-132] ^ d[319-131] ^ d[319-129] ^ d[319-128] ^ d[319-127] ^ d[319-126] ^ d[319-124] ^ d[319-122] ^ d[319-120] ^ d[319-119] ^ d[319-118] ^ d[319-117] ^ d[319-115] ^ d[319-113] ^ d[319-111] ^ d[319-109] ^ d[319-105] ^ d[319-104] ^ d[319-103] ^ d[319-102] ^ d[319-100] ^ d[319-98] ^ d[319-97] ^ d[319-96] ^ d[319-93] ^ d[319-91] ^ d[319-90] ^ d[319-89] ^ d[319-88] ^ d[319-87] ^ d[319-86] ^ d[319-85] ^ d[319-84] ^ d[319-82] ^ d[319-81] ^ d[319-80] ^ d[319-79] ^ d[319-75] ^ d[319-74] ^ d[319-73] ^ d[319-72] ^ d[319-69] ^ d[319-65] ^ d[319-62] ^ d[319-60] ^ d[319-59] ^ d[319-56] ^ d[319-55] ^ d[319-54] ^ d[319-50] ^ d[319-49] ^ d[319-47] ^ d[319-46] ^ d[319-42] ^ d[319-39] ^ d[319-38] ^ d[319-36] ^ d[319-35] ^ d[319-34] ^ d[319-31] ^ d[319-29] ^ d[319-27] ^ d[319-26] ^ d[319-20] ^ d[319-19] ^ d[319-17] ^ d[319-16] ^ d[319-15] ^ d[319-13] ^ d[319-9] ^ d[319-6] ^ d[319-1] ^ d[319-0] ^ c[31-0] ^ c[31-2] ^ c[31-4] ^ c[31-7] ^ c[31-9] ^ c[31-11] ^ c[31-13] ^ c[31-14] ^ c[31-15] ^ c[31-19] ^ c[31-20] ^ c[31-22] ^ c[31-23] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29];
                stage_crc320_crc[7] <= d[319-318] ^ d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-312] ^ d[319-311] ^ d[319-309] ^ d[319-308] ^ d[319-304] ^ d[319-303] ^ d[319-302] ^ d[319-300] ^ d[319-298] ^ d[319-296] ^ d[319-293] ^ d[319-291] ^ d[319-289] ^ d[319-287] ^ d[319-285] ^ d[319-282] ^ d[319-281] ^ d[319-280] ^ d[319-279] ^ d[319-278] ^ d[319-277] ^ d[319-274] ^ d[319-272] ^ d[319-269] ^ d[319-268] ^ d[319-267] ^ d[319-265] ^ d[319-263] ^ d[319-262] ^ d[319-261] ^ d[319-260] ^ d[319-259] ^ d[319-256] ^ d[319-255] ^ d[319-251] ^ d[319-250] ^ d[319-249] ^ d[319-247] ^ d[319-246] ^ d[319-244] ^ d[319-241] ^ d[319-240] ^ d[319-232] ^ d[319-229] ^ d[319-228] ^ d[319-225] ^ d[319-224] ^ d[319-220] ^ d[319-219] ^ d[319-218] ^ d[319-216] ^ d[319-214] ^ d[319-212] ^ d[319-210] ^ d[319-207] ^ d[319-205] ^ d[319-204] ^ d[319-202] ^ d[319-197] ^ d[319-196] ^ d[319-194] ^ d[319-193] ^ d[319-192] ^ d[319-188] ^ d[319-185] ^ d[319-183] ^ d[319-182] ^ d[319-181] ^ d[319-178] ^ d[319-175] ^ d[319-174] ^ d[319-170] ^ d[319-169] ^ d[319-168] ^ d[319-167] ^ d[319-165] ^ d[319-163] ^ d[319-162] ^ d[319-161] ^ d[319-160] ^ d[319-158] ^ d[319-156] ^ d[319-150] ^ d[319-149] ^ d[319-148] ^ d[319-143] ^ d[319-142] ^ d[319-136] ^ d[319-134] ^ d[319-133] ^ d[319-132] ^ d[319-130] ^ d[319-129] ^ d[319-128] ^ d[319-127] ^ d[319-125] ^ d[319-123] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-118] ^ d[319-116] ^ d[319-114] ^ d[319-112] ^ d[319-110] ^ d[319-106] ^ d[319-105] ^ d[319-104] ^ d[319-103] ^ d[319-101] ^ d[319-99] ^ d[319-98] ^ d[319-97] ^ d[319-94] ^ d[319-92] ^ d[319-91] ^ d[319-90] ^ d[319-89] ^ d[319-88] ^ d[319-87] ^ d[319-86] ^ d[319-85] ^ d[319-83] ^ d[319-82] ^ d[319-81] ^ d[319-80] ^ d[319-76] ^ d[319-75] ^ d[319-74] ^ d[319-73] ^ d[319-70] ^ d[319-66] ^ d[319-63] ^ d[319-61] ^ d[319-60] ^ d[319-57] ^ d[319-56] ^ d[319-55] ^ d[319-51] ^ d[319-50] ^ d[319-48] ^ d[319-47] ^ d[319-43] ^ d[319-40] ^ d[319-39] ^ d[319-37] ^ d[319-36] ^ d[319-35] ^ d[319-32] ^ d[319-30] ^ d[319-28] ^ d[319-27] ^ d[319-21] ^ d[319-20] ^ d[319-18] ^ d[319-17] ^ d[319-16] ^ d[319-14] ^ d[319-10] ^ d[319-7] ^ d[319-2] ^ d[319-1] ^ c[31-1] ^ c[31-3] ^ c[31-5] ^ c[31-8] ^ c[31-10] ^ c[31-12] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-20] ^ c[31-21] ^ c[31-23] ^ c[31-24] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30];
                stage_crc320_crc[6] <= d[319-319] ^ d[319-318] ^ d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-313] ^ d[319-312] ^ d[319-310] ^ d[319-309] ^ d[319-305] ^ d[319-304] ^ d[319-303] ^ d[319-301] ^ d[319-299] ^ d[319-297] ^ d[319-294] ^ d[319-292] ^ d[319-290] ^ d[319-288] ^ d[319-286] ^ d[319-283] ^ d[319-282] ^ d[319-281] ^ d[319-280] ^ d[319-279] ^ d[319-278] ^ d[319-275] ^ d[319-273] ^ d[319-270] ^ d[319-269] ^ d[319-268] ^ d[319-266] ^ d[319-264] ^ d[319-263] ^ d[319-262] ^ d[319-261] ^ d[319-260] ^ d[319-257] ^ d[319-256] ^ d[319-252] ^ d[319-251] ^ d[319-250] ^ d[319-248] ^ d[319-247] ^ d[319-245] ^ d[319-242] ^ d[319-241] ^ d[319-233] ^ d[319-230] ^ d[319-229] ^ d[319-226] ^ d[319-225] ^ d[319-221] ^ d[319-220] ^ d[319-219] ^ d[319-217] ^ d[319-215] ^ d[319-213] ^ d[319-211] ^ d[319-208] ^ d[319-206] ^ d[319-205] ^ d[319-203] ^ d[319-198] ^ d[319-197] ^ d[319-195] ^ d[319-194] ^ d[319-193] ^ d[319-189] ^ d[319-186] ^ d[319-184] ^ d[319-183] ^ d[319-182] ^ d[319-179] ^ d[319-176] ^ d[319-175] ^ d[319-171] ^ d[319-170] ^ d[319-169] ^ d[319-168] ^ d[319-166] ^ d[319-164] ^ d[319-163] ^ d[319-162] ^ d[319-161] ^ d[319-159] ^ d[319-157] ^ d[319-151] ^ d[319-150] ^ d[319-149] ^ d[319-144] ^ d[319-143] ^ d[319-137] ^ d[319-135] ^ d[319-134] ^ d[319-133] ^ d[319-131] ^ d[319-130] ^ d[319-129] ^ d[319-128] ^ d[319-126] ^ d[319-124] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-117] ^ d[319-115] ^ d[319-113] ^ d[319-111] ^ d[319-107] ^ d[319-106] ^ d[319-105] ^ d[319-104] ^ d[319-102] ^ d[319-100] ^ d[319-99] ^ d[319-98] ^ d[319-95] ^ d[319-93] ^ d[319-92] ^ d[319-91] ^ d[319-90] ^ d[319-89] ^ d[319-88] ^ d[319-87] ^ d[319-86] ^ d[319-84] ^ d[319-83] ^ d[319-82] ^ d[319-81] ^ d[319-77] ^ d[319-76] ^ d[319-75] ^ d[319-74] ^ d[319-71] ^ d[319-67] ^ d[319-64] ^ d[319-62] ^ d[319-61] ^ d[319-58] ^ d[319-57] ^ d[319-56] ^ d[319-52] ^ d[319-51] ^ d[319-49] ^ d[319-48] ^ d[319-44] ^ d[319-41] ^ d[319-40] ^ d[319-38] ^ d[319-37] ^ d[319-36] ^ d[319-33] ^ d[319-31] ^ d[319-29] ^ d[319-28] ^ d[319-22] ^ d[319-21] ^ d[319-19] ^ d[319-18] ^ d[319-17] ^ d[319-15] ^ d[319-11] ^ d[319-8] ^ d[319-3] ^ d[319-2] ^ c[31-0] ^ c[31-2] ^ c[31-4] ^ c[31-6] ^ c[31-9] ^ c[31-11] ^ c[31-13] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-21] ^ c[31-22] ^ c[31-24] ^ c[31-25] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc320_crc[5] <= d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-313] ^ d[319-312] ^ d[319-311] ^ d[319-309] ^ d[319-306] ^ d[319-304] ^ d[319-303] ^ d[319-299] ^ d[319-297] ^ d[319-296] ^ d[319-294] ^ d[319-293] ^ d[319-292] ^ d[319-291] ^ d[319-290] ^ d[319-289] ^ d[319-288] ^ d[319-286] ^ d[319-284] ^ d[319-282] ^ d[319-281] ^ d[319-280] ^ d[319-277] ^ d[319-273] ^ d[319-271] ^ d[319-270] ^ d[319-268] ^ d[319-267] ^ d[319-263] ^ d[319-262] ^ d[319-259] ^ d[319-258] ^ d[319-255] ^ d[319-253] ^ d[319-251] ^ d[319-249] ^ d[319-246] ^ d[319-242] ^ d[319-237] ^ d[319-231] ^ d[319-228] ^ d[319-224] ^ d[319-222] ^ d[319-221] ^ d[319-220] ^ d[319-218] ^ d[319-210] ^ d[319-208] ^ d[319-206] ^ d[319-204] ^ d[319-203] ^ d[319-202] ^ d[319-201] ^ d[319-197] ^ d[319-196] ^ d[319-195] ^ d[319-193] ^ d[319-192] ^ d[319-191] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-184] ^ d[319-182] ^ d[319-180] ^ d[319-177] ^ d[319-176] ^ d[319-166] ^ d[319-165] ^ d[319-164] ^ d[319-163] ^ d[319-161] ^ d[319-160] ^ d[319-156] ^ d[319-155] ^ d[319-152] ^ d[319-150] ^ d[319-149] ^ d[319-145] ^ d[319-143] ^ d[319-138] ^ d[319-137] ^ d[319-131] ^ d[319-130] ^ d[319-129] ^ d[319-128] ^ d[319-126] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-119] ^ d[319-117] ^ d[319-113] ^ d[319-112] ^ d[319-111] ^ d[319-110] ^ d[319-108] ^ d[319-107] ^ d[319-105] ^ d[319-104] ^ d[319-100] ^ d[319-98] ^ d[319-97] ^ d[319-95] ^ d[319-93] ^ d[319-92] ^ d[319-91] ^ d[319-90] ^ d[319-89] ^ d[319-88] ^ d[319-81] ^ d[319-79] ^ d[319-78] ^ d[319-77] ^ d[319-76] ^ d[319-75] ^ d[319-73] ^ d[319-67] ^ d[319-66] ^ d[319-62] ^ d[319-61] ^ d[319-60] ^ d[319-59] ^ d[319-57] ^ d[319-55] ^ d[319-54] ^ d[319-52] ^ d[319-49] ^ d[319-48] ^ d[319-47] ^ d[319-44] ^ d[319-42] ^ d[319-41] ^ d[319-39] ^ d[319-38] ^ d[319-31] ^ d[319-28] ^ d[319-26] ^ d[319-25] ^ d[319-24] ^ d[319-23] ^ d[319-22] ^ d[319-20] ^ d[319-19] ^ d[319-18] ^ d[319-10] ^ d[319-6] ^ d[319-4] ^ d[319-3] ^ d[319-0] ^ c[31-0] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-8] ^ c[31-9] ^ c[31-11] ^ c[31-15] ^ c[31-16] ^ c[31-18] ^ c[31-21] ^ c[31-23] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28];
                stage_crc320_crc[4] <= d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-313] ^ d[319-312] ^ d[319-310] ^ d[319-307] ^ d[319-305] ^ d[319-304] ^ d[319-300] ^ d[319-298] ^ d[319-297] ^ d[319-295] ^ d[319-294] ^ d[319-293] ^ d[319-292] ^ d[319-291] ^ d[319-290] ^ d[319-289] ^ d[319-287] ^ d[319-285] ^ d[319-283] ^ d[319-282] ^ d[319-281] ^ d[319-278] ^ d[319-274] ^ d[319-272] ^ d[319-271] ^ d[319-269] ^ d[319-268] ^ d[319-264] ^ d[319-263] ^ d[319-260] ^ d[319-259] ^ d[319-256] ^ d[319-254] ^ d[319-252] ^ d[319-250] ^ d[319-247] ^ d[319-243] ^ d[319-238] ^ d[319-232] ^ d[319-229] ^ d[319-225] ^ d[319-223] ^ d[319-222] ^ d[319-221] ^ d[319-219] ^ d[319-211] ^ d[319-209] ^ d[319-207] ^ d[319-205] ^ d[319-204] ^ d[319-203] ^ d[319-202] ^ d[319-198] ^ d[319-197] ^ d[319-196] ^ d[319-194] ^ d[319-193] ^ d[319-192] ^ d[319-189] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-185] ^ d[319-183] ^ d[319-181] ^ d[319-178] ^ d[319-177] ^ d[319-167] ^ d[319-166] ^ d[319-165] ^ d[319-164] ^ d[319-162] ^ d[319-161] ^ d[319-157] ^ d[319-156] ^ d[319-153] ^ d[319-151] ^ d[319-150] ^ d[319-146] ^ d[319-144] ^ d[319-139] ^ d[319-138] ^ d[319-132] ^ d[319-131] ^ d[319-130] ^ d[319-129] ^ d[319-127] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-120] ^ d[319-118] ^ d[319-114] ^ d[319-113] ^ d[319-112] ^ d[319-111] ^ d[319-109] ^ d[319-108] ^ d[319-106] ^ d[319-105] ^ d[319-101] ^ d[319-99] ^ d[319-98] ^ d[319-96] ^ d[319-94] ^ d[319-93] ^ d[319-92] ^ d[319-91] ^ d[319-90] ^ d[319-89] ^ d[319-82] ^ d[319-80] ^ d[319-79] ^ d[319-78] ^ d[319-77] ^ d[319-76] ^ d[319-74] ^ d[319-68] ^ d[319-67] ^ d[319-63] ^ d[319-62] ^ d[319-61] ^ d[319-60] ^ d[319-58] ^ d[319-56] ^ d[319-55] ^ d[319-53] ^ d[319-50] ^ d[319-49] ^ d[319-48] ^ d[319-45] ^ d[319-43] ^ d[319-42] ^ d[319-40] ^ d[319-39] ^ d[319-32] ^ d[319-29] ^ d[319-27] ^ d[319-26] ^ d[319-25] ^ d[319-24] ^ d[319-23] ^ d[319-21] ^ d[319-20] ^ d[319-19] ^ d[319-11] ^ d[319-7] ^ d[319-5] ^ d[319-4] ^ d[319-1] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-9] ^ c[31-10] ^ c[31-12] ^ c[31-16] ^ c[31-17] ^ c[31-19] ^ c[31-22] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29];
                stage_crc320_crc[3] <= d[319-318] ^ d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-313] ^ d[319-311] ^ d[319-308] ^ d[319-306] ^ d[319-305] ^ d[319-301] ^ d[319-299] ^ d[319-298] ^ d[319-296] ^ d[319-295] ^ d[319-294] ^ d[319-293] ^ d[319-292] ^ d[319-291] ^ d[319-290] ^ d[319-288] ^ d[319-286] ^ d[319-284] ^ d[319-283] ^ d[319-282] ^ d[319-279] ^ d[319-275] ^ d[319-273] ^ d[319-272] ^ d[319-270] ^ d[319-269] ^ d[319-265] ^ d[319-264] ^ d[319-261] ^ d[319-260] ^ d[319-257] ^ d[319-255] ^ d[319-253] ^ d[319-251] ^ d[319-248] ^ d[319-244] ^ d[319-239] ^ d[319-233] ^ d[319-230] ^ d[319-226] ^ d[319-224] ^ d[319-223] ^ d[319-222] ^ d[319-220] ^ d[319-212] ^ d[319-210] ^ d[319-208] ^ d[319-206] ^ d[319-205] ^ d[319-204] ^ d[319-203] ^ d[319-199] ^ d[319-198] ^ d[319-197] ^ d[319-195] ^ d[319-194] ^ d[319-193] ^ d[319-190] ^ d[319-189] ^ d[319-188] ^ d[319-187] ^ d[319-186] ^ d[319-184] ^ d[319-182] ^ d[319-179] ^ d[319-178] ^ d[319-168] ^ d[319-167] ^ d[319-166] ^ d[319-165] ^ d[319-163] ^ d[319-162] ^ d[319-158] ^ d[319-157] ^ d[319-154] ^ d[319-152] ^ d[319-151] ^ d[319-147] ^ d[319-145] ^ d[319-140] ^ d[319-139] ^ d[319-133] ^ d[319-132] ^ d[319-131] ^ d[319-130] ^ d[319-128] ^ d[319-124] ^ d[319-123] ^ d[319-122] ^ d[319-121] ^ d[319-119] ^ d[319-115] ^ d[319-114] ^ d[319-113] ^ d[319-112] ^ d[319-110] ^ d[319-109] ^ d[319-107] ^ d[319-106] ^ d[319-102] ^ d[319-100] ^ d[319-99] ^ d[319-97] ^ d[319-95] ^ d[319-94] ^ d[319-93] ^ d[319-92] ^ d[319-91] ^ d[319-90] ^ d[319-83] ^ d[319-81] ^ d[319-80] ^ d[319-79] ^ d[319-78] ^ d[319-77] ^ d[319-75] ^ d[319-69] ^ d[319-68] ^ d[319-64] ^ d[319-63] ^ d[319-62] ^ d[319-61] ^ d[319-59] ^ d[319-57] ^ d[319-56] ^ d[319-54] ^ d[319-51] ^ d[319-50] ^ d[319-49] ^ d[319-46] ^ d[319-44] ^ d[319-43] ^ d[319-41] ^ d[319-40] ^ d[319-33] ^ d[319-30] ^ d[319-28] ^ d[319-27] ^ d[319-26] ^ d[319-25] ^ d[319-24] ^ d[319-22] ^ d[319-21] ^ d[319-20] ^ d[319-12] ^ d[319-8] ^ d[319-6] ^ d[319-5] ^ d[319-2] ^ c[31-0] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-10] ^ c[31-11] ^ c[31-13] ^ c[31-17] ^ c[31-18] ^ c[31-20] ^ c[31-23] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30];
                stage_crc320_crc[2] <= d[319-319] ^ d[319-318] ^ d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-314] ^ d[319-312] ^ d[319-309] ^ d[319-307] ^ d[319-306] ^ d[319-302] ^ d[319-300] ^ d[319-299] ^ d[319-297] ^ d[319-296] ^ d[319-295] ^ d[319-294] ^ d[319-293] ^ d[319-292] ^ d[319-291] ^ d[319-289] ^ d[319-287] ^ d[319-285] ^ d[319-284] ^ d[319-283] ^ d[319-280] ^ d[319-276] ^ d[319-274] ^ d[319-273] ^ d[319-271] ^ d[319-270] ^ d[319-266] ^ d[319-265] ^ d[319-262] ^ d[319-261] ^ d[319-258] ^ d[319-256] ^ d[319-254] ^ d[319-252] ^ d[319-249] ^ d[319-245] ^ d[319-240] ^ d[319-234] ^ d[319-231] ^ d[319-227] ^ d[319-225] ^ d[319-224] ^ d[319-223] ^ d[319-221] ^ d[319-213] ^ d[319-211] ^ d[319-209] ^ d[319-207] ^ d[319-206] ^ d[319-205] ^ d[319-204] ^ d[319-200] ^ d[319-199] ^ d[319-198] ^ d[319-196] ^ d[319-195] ^ d[319-194] ^ d[319-191] ^ d[319-190] ^ d[319-189] ^ d[319-188] ^ d[319-187] ^ d[319-185] ^ d[319-183] ^ d[319-180] ^ d[319-179] ^ d[319-169] ^ d[319-168] ^ d[319-167] ^ d[319-166] ^ d[319-164] ^ d[319-163] ^ d[319-159] ^ d[319-158] ^ d[319-155] ^ d[319-153] ^ d[319-152] ^ d[319-148] ^ d[319-146] ^ d[319-141] ^ d[319-140] ^ d[319-134] ^ d[319-133] ^ d[319-132] ^ d[319-131] ^ d[319-129] ^ d[319-125] ^ d[319-124] ^ d[319-123] ^ d[319-122] ^ d[319-120] ^ d[319-116] ^ d[319-115] ^ d[319-114] ^ d[319-113] ^ d[319-111] ^ d[319-110] ^ d[319-108] ^ d[319-107] ^ d[319-103] ^ d[319-101] ^ d[319-100] ^ d[319-98] ^ d[319-96] ^ d[319-95] ^ d[319-94] ^ d[319-93] ^ d[319-92] ^ d[319-91] ^ d[319-84] ^ d[319-82] ^ d[319-81] ^ d[319-80] ^ d[319-79] ^ d[319-78] ^ d[319-76] ^ d[319-70] ^ d[319-69] ^ d[319-65] ^ d[319-64] ^ d[319-63] ^ d[319-62] ^ d[319-60] ^ d[319-58] ^ d[319-57] ^ d[319-55] ^ d[319-52] ^ d[319-51] ^ d[319-50] ^ d[319-47] ^ d[319-45] ^ d[319-44] ^ d[319-42] ^ d[319-41] ^ d[319-34] ^ d[319-31] ^ d[319-29] ^ d[319-28] ^ d[319-27] ^ d[319-26] ^ d[319-25] ^ d[319-23] ^ d[319-22] ^ d[319-21] ^ d[319-13] ^ d[319-9] ^ d[319-7] ^ d[319-6] ^ d[319-3] ^ c[31-1] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-11] ^ c[31-12] ^ c[31-14] ^ c[31-18] ^ c[31-19] ^ c[31-21] ^ c[31-24] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc320_crc[1] <= d[319-319] ^ d[319-318] ^ d[319-317] ^ d[319-316] ^ d[319-315] ^ d[319-313] ^ d[319-310] ^ d[319-308] ^ d[319-307] ^ d[319-303] ^ d[319-301] ^ d[319-300] ^ d[319-298] ^ d[319-297] ^ d[319-296] ^ d[319-295] ^ d[319-294] ^ d[319-293] ^ d[319-292] ^ d[319-290] ^ d[319-288] ^ d[319-286] ^ d[319-285] ^ d[319-284] ^ d[319-281] ^ d[319-277] ^ d[319-275] ^ d[319-274] ^ d[319-272] ^ d[319-271] ^ d[319-267] ^ d[319-266] ^ d[319-263] ^ d[319-262] ^ d[319-259] ^ d[319-257] ^ d[319-255] ^ d[319-253] ^ d[319-250] ^ d[319-246] ^ d[319-241] ^ d[319-235] ^ d[319-232] ^ d[319-228] ^ d[319-226] ^ d[319-225] ^ d[319-224] ^ d[319-222] ^ d[319-214] ^ d[319-212] ^ d[319-210] ^ d[319-208] ^ d[319-207] ^ d[319-206] ^ d[319-205] ^ d[319-201] ^ d[319-200] ^ d[319-199] ^ d[319-197] ^ d[319-196] ^ d[319-195] ^ d[319-192] ^ d[319-191] ^ d[319-190] ^ d[319-189] ^ d[319-188] ^ d[319-186] ^ d[319-184] ^ d[319-181] ^ d[319-180] ^ d[319-170] ^ d[319-169] ^ d[319-168] ^ d[319-167] ^ d[319-165] ^ d[319-164] ^ d[319-160] ^ d[319-159] ^ d[319-156] ^ d[319-154] ^ d[319-153] ^ d[319-149] ^ d[319-147] ^ d[319-142] ^ d[319-141] ^ d[319-135] ^ d[319-134] ^ d[319-133] ^ d[319-132] ^ d[319-130] ^ d[319-126] ^ d[319-125] ^ d[319-124] ^ d[319-123] ^ d[319-121] ^ d[319-117] ^ d[319-116] ^ d[319-115] ^ d[319-114] ^ d[319-112] ^ d[319-111] ^ d[319-109] ^ d[319-108] ^ d[319-104] ^ d[319-102] ^ d[319-101] ^ d[319-99] ^ d[319-97] ^ d[319-96] ^ d[319-95] ^ d[319-94] ^ d[319-93] ^ d[319-92] ^ d[319-85] ^ d[319-83] ^ d[319-82] ^ d[319-81] ^ d[319-80] ^ d[319-79] ^ d[319-77] ^ d[319-71] ^ d[319-70] ^ d[319-66] ^ d[319-65] ^ d[319-64] ^ d[319-63] ^ d[319-61] ^ d[319-59] ^ d[319-58] ^ d[319-56] ^ d[319-53] ^ d[319-52] ^ d[319-51] ^ d[319-48] ^ d[319-46] ^ d[319-45] ^ d[319-43] ^ d[319-42] ^ d[319-35] ^ d[319-32] ^ d[319-30] ^ d[319-29] ^ d[319-28] ^ d[319-27] ^ d[319-26] ^ d[319-24] ^ d[319-23] ^ d[319-22] ^ d[319-14] ^ d[319-10] ^ d[319-8] ^ d[319-7] ^ d[319-4] ^ c[31-0] ^ c[31-2] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-12] ^ c[31-13] ^ c[31-15] ^ c[31-19] ^ c[31-20] ^ c[31-22] ^ c[31-25] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc320_crc[0] <= d[319-319] ^ d[319-318] ^ d[319-317] ^ d[319-316] ^ d[319-314] ^ d[319-311] ^ d[319-309] ^ d[319-308] ^ d[319-304] ^ d[319-302] ^ d[319-301] ^ d[319-299] ^ d[319-298] ^ d[319-297] ^ d[319-296] ^ d[319-295] ^ d[319-294] ^ d[319-293] ^ d[319-291] ^ d[319-289] ^ d[319-287] ^ d[319-286] ^ d[319-285] ^ d[319-282] ^ d[319-278] ^ d[319-276] ^ d[319-275] ^ d[319-273] ^ d[319-272] ^ d[319-268] ^ d[319-267] ^ d[319-264] ^ d[319-263] ^ d[319-260] ^ d[319-258] ^ d[319-256] ^ d[319-254] ^ d[319-251] ^ d[319-247] ^ d[319-242] ^ d[319-236] ^ d[319-233] ^ d[319-229] ^ d[319-227] ^ d[319-226] ^ d[319-225] ^ d[319-223] ^ d[319-215] ^ d[319-213] ^ d[319-211] ^ d[319-209] ^ d[319-208] ^ d[319-207] ^ d[319-206] ^ d[319-202] ^ d[319-201] ^ d[319-200] ^ d[319-198] ^ d[319-197] ^ d[319-196] ^ d[319-193] ^ d[319-192] ^ d[319-191] ^ d[319-190] ^ d[319-189] ^ d[319-187] ^ d[319-185] ^ d[319-182] ^ d[319-181] ^ d[319-171] ^ d[319-170] ^ d[319-169] ^ d[319-168] ^ d[319-166] ^ d[319-165] ^ d[319-161] ^ d[319-160] ^ d[319-157] ^ d[319-155] ^ d[319-154] ^ d[319-150] ^ d[319-148] ^ d[319-143] ^ d[319-142] ^ d[319-136] ^ d[319-135] ^ d[319-134] ^ d[319-133] ^ d[319-131] ^ d[319-127] ^ d[319-126] ^ d[319-125] ^ d[319-124] ^ d[319-122] ^ d[319-118] ^ d[319-117] ^ d[319-116] ^ d[319-115] ^ d[319-113] ^ d[319-112] ^ d[319-110] ^ d[319-109] ^ d[319-105] ^ d[319-103] ^ d[319-102] ^ d[319-100] ^ d[319-98] ^ d[319-97] ^ d[319-96] ^ d[319-95] ^ d[319-94] ^ d[319-93] ^ d[319-86] ^ d[319-84] ^ d[319-83] ^ d[319-82] ^ d[319-81] ^ d[319-80] ^ d[319-78] ^ d[319-72] ^ d[319-71] ^ d[319-67] ^ d[319-66] ^ d[319-65] ^ d[319-64] ^ d[319-62] ^ d[319-60] ^ d[319-59] ^ d[319-57] ^ d[319-54] ^ d[319-53] ^ d[319-52] ^ d[319-49] ^ d[319-47] ^ d[319-46] ^ d[319-44] ^ d[319-43] ^ d[319-36] ^ d[319-33] ^ d[319-31] ^ d[319-30] ^ d[319-29] ^ d[319-28] ^ d[319-27] ^ d[319-25] ^ d[319-24] ^ d[319-23] ^ d[319-15] ^ d[319-11] ^ d[319-9] ^ d[319-8] ^ d[319-5] ^ c[31-1] ^ c[31-3] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-11] ^ c[31-13] ^ c[31-14] ^ c[31-16] ^ c[31-20] ^ c[31-21] ^ c[31-23] ^ c[31-26] ^ c[31-28] ^ c[31-29] ^ c[31-30] ^ c[31-31];

            end else begin 

                // === CRC32 === 
                
                // Step 0

                // Forward direct signals: valid, last, keep, data_bypass 
                stage_crc32_valid[0] <= stage_masking_valid; 
                stage_crc32_last[0] <= stage_masking_last; 
                stage_crc32_keep[0] <= stage_masking_keep; 
                stage_crc32_data_bypass[0] <= stage_masking_data; 
                stage_crc32_masked_data[0] <= d; 
                crc32_in_flight <= 1'b1; 

                // Reset all other signals of the parallel CRC pipelines 
                stage_crc512_valid <= 1'b0; 
                stage_crc512_last <= 1'b0;
                stage_crc512_keep <= 64'b0; 
                stage_crc512_data_bypass <= 512'b0; 
                stage_crc512_crc <= 32'b0; 

                stage_crc320_valid <= 1'b0; 
                stage_crc320_last <= 1'b0;
                stage_crc320_keep <= 64'b0;
                stage_crc320_data_bypass <= 512'b0; 
                stage_crc320_crc <= 32'b0; 

                // Initialize the valid_stage signal based on the incoming keep 
                if(stage_masking_keep == 64'h000000000000000f) begin 
                    stage_crc32_valid_stages[0][0] <= 1'b1; 
                end else if(stage_masking_keep == 64'h00000000000000ff) begin 
                    stage_crc32_valid_stages[0][1:0] <= 2'b11; 
                end else if(stage_masking_keep == 64'h0000000000000fff) begin
                    stage_crc32_valid_stages[0][2:0] <= 3'b111; 
                end else if(stage_masking_keep == 64'h000000000000ffff) begin 
                    stage_crc32_valid_stages[0][3:0] <= 4'b1111; 
                end

                stage_crc32_crc[0][31] <= d[31-31] ^ d[31-30] ^ d[31-29] ^ d[31-28] ^ d[31-26] ^ d[31-25] ^ d[31-24] ^ d[31-16] ^ d[31-12] ^ d[31-10] ^ d[31-9] ^ d[31-6] ^ d[31-0] ^ c[31-0] ^ c[31-6] ^ c[31-9] ^ c[31-10] ^ c[31-12] ^ c[31-16] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-28] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc32_crc[0][30] <= d[31-28] ^ d[31-27] ^ d[31-24] ^ d[31-17] ^ d[31-16] ^ d[31-13] ^ d[31-12] ^ d[31-11] ^ d[31-9] ^ d[31-7] ^ d[31-6] ^ d[31-1] ^ d[31-0] ^ c[31-0] ^ c[31-1] ^ c[31-6] ^ c[31-7] ^ c[31-9] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-16] ^ c[31-17] ^ c[31-24] ^ c[31-27] ^ c[31-28];
                stage_crc32_crc[0][29] <= d[31-31] ^ d[31-30] ^ d[31-26] ^ d[31-24] ^ d[31-18] ^ d[31-17] ^ d[31-16] ^ d[31-14] ^ d[31-13] ^ d[31-9] ^ d[31-8] ^ d[31-7] ^ d[31-6] ^ d[31-2] ^ d[31-1] ^ d[31-0] ^ c[31-0] ^ c[31-1] ^ c[31-2] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-13] ^ c[31-14] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-24] ^ c[31-26] ^ c[31-30] ^ c[31-31];
                stage_crc32_crc[0][28] <= d[31-31] ^ d[31-27] ^ d[31-25] ^ d[31-19] ^ d[31-18] ^ d[31-17] ^ d[31-15] ^ d[31-14] ^ d[31-10] ^ d[31-9] ^ d[31-8] ^ d[31-7] ^ d[31-3] ^ d[31-2] ^ d[31-1] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-10] ^ c[31-14] ^ c[31-15] ^ c[31-17] ^ c[31-18] ^ c[31-19] ^ c[31-25] ^ c[31-27] ^ c[31-31];
                stage_crc32_crc[0][27] <= d[31-31] ^ d[31-30] ^ d[31-29] ^ d[31-25] ^ d[31-24] ^ d[31-20] ^ d[31-19] ^ d[31-18] ^ d[31-15] ^ d[31-12] ^ d[31-11] ^ d[31-8] ^ d[31-6] ^ d[31-4] ^ d[31-3] ^ d[31-2] ^ d[31-0] ^ c[31-0] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-6] ^ c[31-8] ^ c[31-11] ^ c[31-12] ^ c[31-15] ^ c[31-18] ^ c[31-19] ^ c[31-20] ^ c[31-24] ^ c[31-25] ^ c[31-29] ^ c[31-30] ^ c[31-31];
                stage_crc32_crc[0][26] <= d[31-29] ^ d[31-28] ^ d[31-24] ^ d[31-21] ^ d[31-20] ^ d[31-19] ^ d[31-13] ^ d[31-10] ^ d[31-7] ^ d[31-6] ^ d[31-5] ^ d[31-4] ^ d[31-3] ^ d[31-1] ^ d[31-0] ^ c[31-0] ^ c[31-1] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-10] ^ c[31-13] ^ c[31-19] ^ c[31-20] ^ c[31-21] ^ c[31-24] ^ c[31-28] ^ c[31-29];
                stage_crc32_crc[0][25] <= d[31-30] ^ d[31-29] ^ d[31-25] ^ d[31-22] ^ d[31-21] ^ d[31-20] ^ d[31-14] ^ d[31-11] ^ d[31-8] ^ d[31-7] ^ d[31-6] ^ d[31-5] ^ d[31-4] ^ d[31-2] ^ d[31-1] ^ c[31-1] ^ c[31-2] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-11] ^ c[31-14] ^ c[31-20] ^ c[31-21] ^ c[31-22] ^ c[31-25] ^ c[31-29] ^ c[31-30];
                stage_crc32_crc[0][24] <= d[31-29] ^ d[31-28] ^ d[31-25] ^ d[31-24] ^ d[31-23] ^ d[31-22] ^ d[31-21] ^ d[31-16] ^ d[31-15] ^ d[31-10] ^ d[31-8] ^ d[31-7] ^ d[31-5] ^ d[31-3] ^ d[31-2] ^ d[31-0] ^ c[31-0] ^ c[31-2] ^ c[31-3] ^ c[31-5] ^ c[31-7] ^ c[31-8] ^ c[31-10] ^ c[31-15] ^ c[31-16] ^ c[31-21] ^ c[31-22] ^ c[31-23] ^ c[31-24] ^ c[31-25] ^ c[31-28] ^ c[31-29];
                stage_crc32_crc[0][23] <= d[31-31] ^ d[31-28] ^ d[31-23] ^ d[31-22] ^ d[31-17] ^ d[31-12] ^ d[31-11] ^ d[31-10] ^ d[31-8] ^ d[31-4] ^ d[31-3] ^ d[31-1] ^ d[31-0] ^ c[31-0] ^ c[31-1] ^ c[31-3] ^ c[31-4] ^ c[31-8] ^ c[31-10] ^ c[31-11] ^ c[31-12] ^ c[31-17] ^ c[31-22] ^ c[31-23] ^ c[31-28] ^ c[31-31];
                stage_crc32_crc[0][22] <= d[31-29] ^ d[31-24] ^ d[31-23] ^ d[31-18] ^ d[31-13] ^ d[31-12] ^ d[31-11] ^ d[31-9] ^ d[31-5] ^ d[31-4] ^ d[31-2] ^ d[31-1] ^ c[31-1] ^ c[31-2] ^ c[31-4] ^ c[31-5] ^ c[31-9] ^ c[31-11] ^ c[31-12] ^ c[31-13] ^ c[31-18] ^ c[31-23] ^ c[31-24] ^ c[31-29];
                stage_crc32_crc[0][21] <= d[31-31] ^ d[31-29] ^ d[31-28] ^ d[31-26] ^ d[31-19] ^ d[31-16] ^ d[31-14] ^ d[31-13] ^ d[31-9] ^ d[31-5] ^ d[31-3] ^ d[31-2] ^ d[31-0] ^ c[31-0] ^ c[31-2] ^ c[31-3] ^ c[31-5] ^ c[31-9] ^ c[31-13] ^ c[31-14] ^ c[31-16] ^ c[31-19] ^ c[31-26] ^ c[31-28] ^ c[31-29] ^ c[31-31];
                stage_crc32_crc[0][20] <= d[31-31] ^ d[31-28] ^ d[31-27] ^ d[31-26] ^ d[31-25] ^ d[31-24] ^ d[31-20] ^ d[31-17] ^ d[31-16] ^ d[31-15] ^ d[31-14] ^ d[31-12] ^ d[31-9] ^ d[31-4] ^ d[31-3] ^ d[31-1] ^ d[31-0] ^ c[31-0] ^ c[31-1] ^ c[31-3] ^ c[31-4] ^ c[31-9] ^ c[31-12] ^ c[31-14] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-20] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-31];
                stage_crc32_crc[0][19] <= d[31-31] ^ d[31-30] ^ d[31-27] ^ d[31-24] ^ d[31-21] ^ d[31-18] ^ d[31-17] ^ d[31-15] ^ d[31-13] ^ d[31-12] ^ d[31-9] ^ d[31-6] ^ d[31-5] ^ d[31-4] ^ d[31-2] ^ d[31-1] ^ d[31-0] ^ c[31-0] ^ c[31-1] ^ c[31-2] ^ c[31-4] ^ c[31-5] ^ c[31-6] ^ c[31-9] ^ c[31-12] ^ c[31-13] ^ c[31-15] ^ c[31-17] ^ c[31-18] ^ c[31-21] ^ c[31-24] ^ c[31-27] ^ c[31-30] ^ c[31-31];
                stage_crc32_crc[0][18] <= d[31-31] ^ d[31-28] ^ d[31-25] ^ d[31-22] ^ d[31-19] ^ d[31-18] ^ d[31-16] ^ d[31-14] ^ d[31-13] ^ d[31-10] ^ d[31-7] ^ d[31-6] ^ d[31-5] ^ d[31-3] ^ d[31-2] ^ d[31-1] ^ c[31-1] ^ c[31-2] ^ c[31-3] ^ c[31-5] ^ c[31-6] ^ c[31-7] ^ c[31-10] ^ c[31-13] ^ c[31-14] ^ c[31-16] ^ c[31-18] ^ c[31-19] ^ c[31-22] ^ c[31-25] ^ c[31-28] ^ c[31-31];
                stage_crc32_crc[0][17] <= d[31-29] ^ d[31-26] ^ d[31-23] ^ d[31-20] ^ d[31-19] ^ d[31-17] ^ d[31-15] ^ d[31-14] ^ d[31-11] ^ d[31-8] ^ d[31-7] ^ d[31-6] ^ d[31-4] ^ d[31-3] ^ d[31-2] ^ c[31-2] ^ c[31-3] ^ c[31-4] ^ c[31-6] ^ c[31-7] ^ c[31-8] ^ c[31-11] ^ c[31-14] ^ c[31-15] ^ c[31-17] ^ c[31-19] ^ c[31-20] ^ c[31-23] ^ c[31-26] ^ c[31-29];
                stage_crc32_crc[0][16] <= d[31-30] ^ d[31-27] ^ d[31-24] ^ d[31-21] ^ d[31-20] ^ d[31-18] ^ d[31-16] ^ d[31-15] ^ d[31-12] ^ d[31-9] ^ d[31-8] ^ d[31-7] ^ d[31-5] ^ d[31-4] ^ d[31-3] ^ c[31-3] ^ c[31-4] ^ c[31-5] ^ c[31-7] ^ c[31-8] ^ c[31-9] ^ c[31-12] ^ c[31-15] ^ c[31-16] ^ c[31-18] ^ c[31-20] ^ c[31-21] ^ c[31-24] ^ c[31-27] ^ c[31-30];
                stage_crc32_crc[0][15] <= d[31-30] ^ d[31-29] ^ d[31-26] ^ d[31-24] ^ d[31-22] ^ d[31-21] ^ d[31-19] ^ d[31-17] ^ d[31-13] ^ d[31-12] ^ d[31-8] ^ d[31-5] ^ d[31-4] ^ d[31-0] ^ c[31-0] ^ c[31-4] ^ c[31-5] ^ c[31-8] ^ c[31-12] ^ c[31-13] ^ c[31-17] ^ c[31-19] ^ c[31-21] ^ c[31-22] ^ c[31-24] ^ c[31-26] ^ c[31-29] ^ c[31-30];
                stage_crc32_crc[0][14] <= d[31-31] ^ d[31-30] ^ d[31-27] ^ d[31-25] ^ d[31-23] ^ d[31-22] ^ d[31-20] ^ d[31-18] ^ d[31-14] ^ d[31-13] ^ d[31-9] ^ d[31-6] ^ d[31-5] ^ d[31-1] ^ c[31-1] ^ c[31-5] ^ c[31-6] ^ c[31-9] ^ c[31-13] ^ c[31-14] ^ c[31-18] ^ c[31-20] ^ c[31-22] ^ c[31-23] ^ c[31-25] ^ c[31-27] ^ c[31-30] ^ c[31-31];
                stage_crc32_crc[0][13] <= d[31-31] ^ d[31-28] ^ d[31-26] ^ d[31-24] ^ d[31-23] ^ d[31-21] ^ d[31-19] ^ d[31-15] ^ d[31-14] ^ d[31-10] ^ d[31-7] ^ d[31-6] ^ d[31-2] ^ c[31-2] ^ c[31-6] ^ c[31-7] ^ c[31-10] ^ c[31-14] ^ c[31-15] ^ c[31-19] ^ c[31-21] ^ c[31-23] ^ c[31-24] ^ c[31-26] ^ c[31-28] ^ c[31-31];
                stage_crc32_crc[0][12] <= d[31-29] ^ d[31-27] ^ d[31-25] ^ d[31-24] ^ d[31-22] ^ d[31-20] ^ d[31-16] ^ d[31-15] ^ d[31-11] ^ d[31-8] ^ d[31-7] ^ d[31-3] ^ c[31-3] ^ c[31-7] ^ c[31-8] ^ c[31-11] ^ c[31-15] ^ c[31-16] ^ c[31-20] ^ c[31-22] ^ c[31-24] ^ c[31-25] ^ c[31-27] ^ c[31-29];
                stage_crc32_crc[0][11] <= d[31-30] ^ d[31-28] ^ d[31-26] ^ d[31-25] ^ d[31-23] ^ d[31-21] ^ d[31-17] ^ d[31-16] ^ d[31-12] ^ d[31-9] ^ d[31-8] ^ d[31-4] ^ c[31-4] ^ c[31-8] ^ c[31-9] ^ c[31-12] ^ c[31-16] ^ c[31-17] ^ c[31-21] ^ c[31-23] ^ c[31-25] ^ c[31-26] ^ c[31-28] ^ c[31-30];
                stage_crc32_crc[0][10] <= d[31-31] ^ d[31-29] ^ d[31-27] ^ d[31-26] ^ d[31-24] ^ d[31-22] ^ d[31-18] ^ d[31-17] ^ d[31-13] ^ d[31-10] ^ d[31-9] ^ d[31-5] ^ c[31-5] ^ c[31-9] ^ c[31-10] ^ c[31-13] ^ c[31-17] ^ c[31-18] ^ c[31-22] ^ c[31-24] ^ c[31-26] ^ c[31-27] ^ c[31-29] ^ c[31-31];
                stage_crc32_crc[0][9] <= d[31-31] ^ d[31-29] ^ d[31-27] ^ d[31-26] ^ d[31-24] ^ d[31-23] ^ d[31-19] ^ d[31-18] ^ d[31-16] ^ d[31-14] ^ d[31-12] ^ d[31-11] ^ d[31-9] ^ d[31-0] ^ c[31-0] ^ c[31-9] ^ c[31-11] ^ c[31-12] ^ c[31-14] ^ c[31-16] ^ c[31-18] ^ c[31-19] ^ c[31-23] ^ c[31-24] ^ c[31-26] ^ c[31-27] ^ c[31-29] ^ c[31-31];
                stage_crc32_crc[0][8] <= d[31-31] ^ d[31-29] ^ d[31-27] ^ d[31-26] ^ d[31-20] ^ d[31-19] ^ d[31-17] ^ d[31-16] ^ d[31-15] ^ d[31-13] ^ d[31-9] ^ d[31-6] ^ d[31-1] ^ d[31-0] ^ c[31-0] ^ c[31-1] ^ c[31-6] ^ c[31-9] ^ c[31-13] ^ c[31-15] ^ c[31-16] ^ c[31-17] ^ c[31-19] ^ c[31-20] ^ c[31-26] ^ c[31-27] ^ c[31-29] ^ c[31-31];
                stage_crc32_crc[0][7] <= d[31-30] ^ d[31-28] ^ d[31-27] ^ d[31-21] ^ d[31-20] ^ d[31-18] ^ d[31-17] ^ d[31-16] ^ d[31-14] ^ d[31-10] ^ d[31-7] ^ d[31-2] ^ d[31-1] ^ c[31-1] ^ c[31-2] ^ c[31-7] ^ c[31-10] ^ c[31-14] ^ c[31-16] ^ c[31-17] ^ c[31-18] ^ c[31-20] ^ c[31-21] ^ c[31-27] ^ c[31-28] ^ c[31-30];
                stage_crc32_crc[0][6] <= d[31-31] ^ d[31-29] ^ d[31-28] ^ d[31-22] ^ d[31-21] ^ d[31-19] ^ d[31-18] ^ d[31-17] ^ d[31-15] ^ d[31-11] ^ d[31-8] ^ d[31-3] ^ d[31-2] ^ c[31-2] ^ c[31-3] ^ c[31-8] ^ c[31-11] ^ c[31-15] ^ c[31-17] ^ c[31-18] ^ c[31-19] ^ c[31-21] ^ c[31-22] ^ c[31-28] ^ c[31-29] ^ c[31-31];
                stage_crc32_crc[0][5] <= d[31-31] ^ d[31-28] ^ d[31-26] ^ d[31-25] ^ d[31-24] ^ d[31-23] ^ d[31-22] ^ d[31-20] ^ d[31-19] ^ d[31-18] ^ d[31-10] ^ d[31-6] ^ d[31-4] ^ d[31-3] ^ d[31-0] ^ c[31-0] ^ c[31-3] ^ c[31-4] ^ c[31-6] ^ c[31-10] ^ c[31-18] ^ c[31-19] ^ c[31-20] ^ c[31-22] ^ c[31-23] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-28] ^ c[31-31];
                stage_crc32_crc[0][4] <= d[31-29] ^ d[31-27] ^ d[31-26] ^ d[31-25] ^ d[31-24] ^ d[31-23] ^ d[31-21] ^ d[31-20] ^ d[31-19] ^ d[31-11] ^ d[31-7] ^ d[31-5] ^ d[31-4] ^ d[31-1] ^ c[31-1] ^ c[31-4] ^ c[31-5] ^ c[31-7] ^ c[31-11] ^ c[31-19] ^ c[31-20] ^ c[31-21] ^ c[31-23] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-29];
                stage_crc32_crc[0][3] <= d[31-30] ^ d[31-28] ^ d[31-27] ^ d[31-26] ^ d[31-25] ^ d[31-24] ^ d[31-22] ^ d[31-21] ^ d[31-20] ^ d[31-12] ^ d[31-8] ^ d[31-6] ^ d[31-5] ^ d[31-2] ^ c[31-2] ^ c[31-5] ^ c[31-6] ^ c[31-8] ^ c[31-12] ^ c[31-20] ^ c[31-21] ^ c[31-22] ^ c[31-24] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-30];
                stage_crc32_crc[0][2] <= d[31-31] ^ d[31-29] ^ d[31-28] ^ d[31-27] ^ d[31-26] ^ d[31-25] ^ d[31-23] ^ d[31-22] ^ d[31-21] ^ d[31-13] ^ d[31-9] ^ d[31-7] ^ d[31-6] ^ d[31-3] ^ c[31-3] ^ c[31-6] ^ c[31-7] ^ c[31-9] ^ c[31-13] ^ c[31-21] ^ c[31-22] ^ c[31-23] ^ c[31-25] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-31];
                stage_crc32_crc[0][1] <= d[31-30] ^ d[31-29] ^ d[31-28] ^ d[31-27] ^ d[31-26] ^ d[31-24] ^ d[31-23] ^ d[31-22] ^ d[31-14] ^ d[31-10] ^ d[31-8] ^ d[31-7] ^ d[31-4] ^ c[31-4] ^ c[31-7] ^ c[31-8] ^ c[31-10] ^ c[31-14] ^ c[31-22] ^ c[31-23] ^ c[31-24] ^ c[31-26] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30];
                stage_crc32_crc[0][0] <= d[31-31] ^ d[31-30] ^ d[31-29] ^ d[31-28] ^ d[31-27] ^ d[31-25] ^ d[31-24] ^ d[31-23] ^ d[31-15] ^ d[31-11] ^ d[31-9] ^ d[31-8] ^ d[31-5] ^ c[31-5] ^ c[31-8] ^ c[31-9] ^ c[31-11] ^ c[31-15] ^ c[31-23] ^ c[31-24] ^ c[31-25] ^ c[31-27] ^ c[31-28] ^ c[31-29] ^ c[31-30] ^ c[31-31];


                // // Step 1 - 15, written down in a parallelized for-loop 
                // for(integer stage = 1; stage < 16; stage++) begin

                //     // Forward direct signals: valid, last, keep, data_bypass 
                //     stage_crc32_valid[stage] <= stage_crc32_valid[stage-1];
                //     stage_crc32_last[stage] <= stage_crc32_last[stage-1]; 
                //     stage_crc32_keep[stage] <= stage_crc32_keep[stage-1]; 
                //     stage_crc32_data_bypass[stage] <= stage_crc32_data_bypass[stage-1]; 
                //     stage_crc32_masked_data[stage] <= stage_crc32_masked_data[stage-1]; 

                //     // Calculate the CRC-value if the keep signal indicates that the part of the dataword is still valid 
                //     if(stage_crc32_keep_stage[stage] == 4'hf) begin 
                //         crc32_test_probe <= 1'b1; 

                //         stage_crc32_crc[stage][31] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][30] <= stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28];
                //         stage_crc32_crc[stage][29] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][28] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][27] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][26] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29];
                //         stage_crc32_crc[stage][25] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30];
                //         stage_crc32_crc[stage][24] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29];
                //         stage_crc32_crc[stage][23] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][22] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-29];
                //         stage_crc32_crc[stage][21] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][20] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][19] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][18] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][17] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-29];
                //         stage_crc32_crc[stage][16] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-30];
                //         stage_crc32_crc[stage][15] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30];
                //         stage_crc32_crc[stage][14] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][13] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][12] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29];
                //         stage_crc32_crc[stage][11] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-30];
                //         stage_crc32_crc[stage][10] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][9] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][8] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][7] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-30];
                //         stage_crc32_crc[stage][6] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][5] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][4] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29];
                //         stage_crc32_crc[stage][3] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-30];
                //         stage_crc32_crc[stage][2] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                //         stage_crc32_crc[stage][1] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30];
                //         stage_crc32_crc[stage][0] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];

                //     end else begin 
                //         stage_crc32_crc[stage] <= stage_crc32_crc[stage-1];  
                //     end 
                // end 

            end 

        end else begin 
            // If previous stage is not valid anymore, all signals in the CRC-stage should be reset 
            stage_crc512_valid <= 1'b0; 
            stage_crc512_last <= 1'b0; 
            stage_crc512_keep <= 64'b0; 
            stage_crc512_data_bypass <= 512'b0; 

            if(!stage_crc_follow_up_word) begin 
                stage_crc512_crc <= 32'b0;
            end

            stage_crc320_valid <= 1'b0; 
            stage_crc320_last <= 1'b0; 
            stage_crc320_keep <= 64'b0; 
            stage_crc320_data_bypass <= 512'b0; 
            stage_crc320_crc <= 32'b0; 

            stage_crc32_valid[0] <= 1'b0; 
            stage_crc32_last[0] <= 1'b0; 
            stage_crc32_keep[0] <= 64'b0; 
            stage_crc32_data_bypass[0] <= 512'b0; 
            stage_crc32_masked_data[0] <= 512'b0; 
            stage_crc32_crc[0] <= 32'b0; 

        end 


        ///////////////////////////////////////////////////////////////////////
        //
        // STAGE(S) 2.5: REST OF THE CRC32-PIPELINE
        //
        ///////////////////////////////////////////////////////////////////////

        for(integer stage = 1; stage < 16; stage++) begin
            if(!stage_crc32_early_done) begin 
                stage_crc32_valid[stage] <= stage_crc32_valid[stage-1]; 
                stage_crc32_last[stage] <= stage_crc32_last[stage-1];
                stage_crc32_keep[stage] <= stage_crc32_keep[stage-1]; 
                stage_crc32_data_bypass[stage] <= stage_crc32_data_bypass[stage-1]; 
                stage_crc32_masked_data[stage] <= stage_crc32_masked_data[stage-1]; 
            end else begin 
                stage_crc32_valid[stage] <= 1'b0; 
                stage_crc32_last[stage] <= 1'b0; 
                stage_crc32_keep[stage] <= 64'b0;
                stage_crc32_data_bypass[stage] <= 512'b0;
                stage_crc32_masked_data[stage] <= 512'b0; 
            end 

            if(stage_crc32_valid[stage-1]) begin 
                // Calculate the CRC-value if the keep signal indicates that the part of the dataword is still valid 
                if(stage_crc32_keep_stage[stage] == 4'hf) begin 
                    crc32_test_probe <= 1'b1; 

                    stage_crc32_crc[stage][31] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][30] <= stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28];
                    stage_crc32_crc[stage][29] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][28] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][27] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][26] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29];
                    stage_crc32_crc[stage][25] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30];
                    stage_crc32_crc[stage][24] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29];
                    stage_crc32_crc[stage][23] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][22] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-29];
                    stage_crc32_crc[stage][21] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][20] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][19] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][18] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][17] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-29];
                    stage_crc32_crc[stage][16] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-30];
                    stage_crc32_crc[stage][15] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30];
                    stage_crc32_crc[stage][14] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][13] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][12] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29];
                    stage_crc32_crc[stage][11] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-30];
                    stage_crc32_crc[stage][10] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][9] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][8] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][7] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-16+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-16] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-30];
                    stage_crc32_crc[stage][6] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-17+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-17] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][5] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-18+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_masked_data[stage-1][31-0+stage*32] ^ stage_crc32_crc[stage-1][31-0] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-18] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][4] <= stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-19+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_masked_data[stage-1][31-1+stage*32] ^ stage_crc32_crc[stage-1][31-1] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-19] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-29];
                    stage_crc32_crc[stage][3] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-20+stage*32] ^ stage_crc32_masked_data[stage-1][31-12+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_masked_data[stage-1][31-2+stage*32] ^ stage_crc32_crc[stage-1][31-2] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-12] ^ stage_crc32_crc[stage-1][31-20] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-30];
                    stage_crc32_crc[stage][2] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-21+stage*32] ^ stage_crc32_masked_data[stage-1][31-13+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-6+stage*32] ^ stage_crc32_masked_data[stage-1][31-3+stage*32] ^ stage_crc32_crc[stage-1][31-3] ^ stage_crc32_crc[stage-1][31-6] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-13] ^ stage_crc32_crc[stage-1][31-21] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-31];
                    stage_crc32_crc[stage][1] <= stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-26+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-22+stage*32] ^ stage_crc32_masked_data[stage-1][31-14+stage*32] ^ stage_crc32_masked_data[stage-1][31-10+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-7+stage*32] ^ stage_crc32_masked_data[stage-1][31-4+stage*32] ^ stage_crc32_crc[stage-1][31-4] ^ stage_crc32_crc[stage-1][31-7] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-10] ^ stage_crc32_crc[stage-1][31-14] ^ stage_crc32_crc[stage-1][31-22] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-26] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30];
                    stage_crc32_crc[stage][0] <= stage_crc32_masked_data[stage-1][31-31+stage*32] ^ stage_crc32_masked_data[stage-1][31-30+stage*32] ^ stage_crc32_masked_data[stage-1][31-29+stage*32] ^ stage_crc32_masked_data[stage-1][31-28+stage*32] ^ stage_crc32_masked_data[stage-1][31-27+stage*32] ^ stage_crc32_masked_data[stage-1][31-25+stage*32] ^ stage_crc32_masked_data[stage-1][31-24+stage*32] ^ stage_crc32_masked_data[stage-1][31-23+stage*32] ^ stage_crc32_masked_data[stage-1][31-15+stage*32] ^ stage_crc32_masked_data[stage-1][31-11+stage*32] ^ stage_crc32_masked_data[stage-1][31-9+stage*32] ^ stage_crc32_masked_data[stage-1][31-8+stage*32] ^ stage_crc32_masked_data[stage-1][31-5+stage*32] ^ stage_crc32_crc[stage-1][31-5] ^ stage_crc32_crc[stage-1][31-8] ^ stage_crc32_crc[stage-1][31-9] ^ stage_crc32_crc[stage-1][31-11] ^ stage_crc32_crc[stage-1][31-15] ^ stage_crc32_crc[stage-1][31-23] ^ stage_crc32_crc[stage-1][31-24] ^ stage_crc32_crc[stage-1][31-25] ^ stage_crc32_crc[stage-1][31-27] ^ stage_crc32_crc[stage-1][31-28] ^ stage_crc32_crc[stage-1][31-29] ^ stage_crc32_crc[stage-1][31-30] ^ stage_crc32_crc[stage-1][31-31];

                end else begin 
                    stage_crc32_crc[stage] <= stage_crc32_crc[stage-1];  
                    if(!stage_crc32_early_done) begin 
                        stage_crc32_early_done <= 1'b1; 
                        stage_crc32_counter_word <= stage; 
                    end 
                end 
            end else begin
                stage_crc32_crc[stage] <= 32'b0; 
            end 
        end

        ///////////////////////////////////////////////////////////////////////
        //
        // STAGE 3: JOIN CRC-PIPELINES
        //
        ////////////////////////////////////////////////////////////////////////

        // Find out which of the three CRC-pipelines is firing at the moment and adopt its value 
        if(stage_crc512_valid) begin 
            stage_join_valid <= stage_crc512_valid; 
            stage_join_data <= stage_crc512_data_bypass; 
            stage_join_crc <= stage_crc512_crc ^ 32'hffffffff; 
            stage_join_keep <= stage_crc512_keep; 
            stage_join_last <= stage_crc512_last; 
        end else if(stage_crc320_valid) begin 
            stage_join_valid <= stage_crc320_valid; 
            stage_join_data <= stage_crc320_data_bypass; 
            stage_join_crc <= stage_crc320_crc ^ 32'hffffffff; 
            stage_join_keep <= stage_crc320_keep; 
            stage_join_last <= stage_crc320_last; 
        end else if(stage_crc32_valid[15]) begin 
            stage_join_valid <= stage_crc32_valid[15];
            stage_join_data <= stage_crc32_data_bypass[15]; 
            stage_join_crc <= stage_crc32_crc[15] ^ 32'hffffffff; 
            stage_join_keep <= stage_crc32_keep[15]; 
            stage_join_last <= stage_crc32_last[15]; 
            crc32_in_flight <= 1'b0; 
        end else if(stage_crc32_early_done) begin
            stage_join_valid <= stage_crc32_valid[stage_crc32_counter_word]; 
            stage_join_crc <= stage_crc32_crc[stage_crc32_counter_word] ^32'hffffffff; 
            stage_join_data <= stage_crc32_data_bypass[stage_crc32_counter_word]; 
            stage_join_keep <= stage_crc32_keep[stage_crc32_counter_word];
            stage_join_last <= stage_crc32_last[stage_crc32_counter_word]; 
            stage_crc32_early_done <= 0;
            stage_crc32_counter_word <= 4'b0; 
            crc32_in_flight <= 1'b0; 
        end else begin 
            stage_join_valid <= 1'b0; 
            stage_join_data <= 512'b0; 
            stage_join_crc <= 32'b0; 
            stage_join_keep <= 64'b0; 
            stage_join_last <= 1'b0; 
        end


        ///////////////////////////////////////////////////////////////////////
        //
        // STAGE 4: CRC INSERTION
        //
        ///////////////////////////////////////////////////////////////////////
        
        // If not last, value must be forwarded without crc-insertion to be picked up at output
        if(!stage_join_last) begin 
            // Forward direct values: valid, last, keep 
            stage_reinsertion_valid <= stage_join_valid; 
            stage_reinsertion_last <= stage_join_last; 
            stage_reinsertion_keep <= stage_join_keep; 
            stage_reinsertion_data <= stage_join_data; 
            stage_reinsertion_crc <= stage_join_crc; 

        // If the word is last, previously calculated CRC-value needs to be inserted before the word can be picked up at output    
        end else begin 
            // Pass on valid anyways 
            stage_reinsertion_valid <= stage_join_valid; 

            // Based on keep, check if the word is full 
            if(stage_join_keep[63] == 1'b1) begin
                stage_reinsertion_last <= 0; 
                stage_reinsertion_data <= stage_join_data;
                stage_reinsertion_crc <= stage_join_crc; 
                stage_reinsertion_keep <= stage_join_keep;

                // In this case, the pipeline must be stalled for one cycle to include the freshly formed word 
                stall_pipeline <= 1'b1; 

            end else begin 
                // Pass on last 
                stage_reinsertion_last <= stage_join_last; 
                stall_pipeline <= 1'b0; 

                if(stage_join_keep == 4'hf) begin
                    stage_reinsertion_data[31:0] <= stage_join_data[31:0];
                    stage_reinsertion_data[63:32] <= stage_join_crc; 
                    stage_reinsertion_data[511:64] <= 448'b0; 
                    stage_reinsertion_keep[7:0] <= 8'hff;
                    stage_reinsertion_keep[63:8] <= 56'h0;
                end else if(stage_join_keep == 8'hff) begin 
                    stage_reinsertion_data[63:0] <= stage_join_data[63:0]; 
                    stage_reinsertion_data[95:64] <= stage_join_crc; 
                    stage_reinsertion_data[511:96] <= 416'b0; 
                    stage_reinsertion_keep[11:0] <= 12'hfff;
                    stage_reinsertion_keep[63:12] <= 52'h0;
                end else if(stage_join_keep == 12'hfff) begin 
                    stage_reinsertion_data[95:0] <= stage_join_data[95:0]; 
                    stage_reinsertion_data[127:96] <= stage_join_crc; 
                    stage_reinsertion_data[511:128] <= 384'b0; 
                    stage_reinsertion_keep[15:0] <= 16'hffff;
                    stage_reinsertion_keep[63:16] <= 48'h0;
                end else if(stage_join_keep == 16'hffff) begin 
                    stage_reinsertion_data[127:0] <= stage_join_data[127:0]; 
                    stage_reinsertion_data[159:128] <= stage_join_crc; 
                    stage_reinsertion_data[511:160] <= 352'b0; 
                    stage_reinsertion_keep[19:0] <= 20'hfffff;
                    stage_reinsertion_keep[63:20] <= 44'h0;
                end else if(stage_join_keep == 20'hfffff) begin 
                    stage_reinsertion_data[159:0] <= stage_join_data[159:0]; 
                    stage_reinsertion_data[191:160] <= stage_join_crc; 
                    stage_reinsertion_data[511:192] <= 320'b0; 
                    stage_reinsertion_keep[23:0] <= 24'hffffff;
                    stage_reinsertion_keep[63:24] <= 40'h0;
                end else if(stage_join_keep == 24'hffffff) begin 
                    stage_reinsertion_data[191:0] <= stage_join_data[191:0]; 
                    stage_reinsertion_data[223:192] <= stage_join_crc; 
                    stage_reinsertion_data[511:224] <= 288'b0; 
                    stage_reinsertion_keep[27:0] <= 28'hfffffff;
                    stage_reinsertion_keep[63:28] <= 36'h0;
                end else if(stage_join_keep == 28'hfffffff) begin
                    stage_reinsertion_data[223:0] <= stage_join_data[223:0]; 
                    stage_reinsertion_data[255:224] <= stage_join_crc; 
                    stage_reinsertion_data[511:256] <= 256'b0; 
                    stage_reinsertion_keep[31:0] <= 32'hffffffff;
                    stage_reinsertion_keep[63:32] <= 32'h0;
                end else if(stage_join_keep == 32'hffffffff) begin 
                    stage_reinsertion_data[255:0] <= stage_join_data[255:0]; 
                    stage_reinsertion_data[287:256] <= stage_join_crc; 
                    stage_reinsertion_data[511:288] <= 224'b0; 
                    stage_reinsertion_keep[35:0] <= 36'hfffffffff;
                    stage_reinsertion_keep[63:36] <= 28'h0;
                end else if(stage_join_keep == 36'hfffffffff) begin
                    stage_reinsertion_data[287:0] <= stage_join_data[287:0]; 
                    stage_reinsertion_data[319:288] <= stage_join_crc; 
                    stage_reinsertion_data[511:320] <= 192'b0; 
                    stage_reinsertion_keep[39:0] <= 40'hffffffffff;
                    stage_reinsertion_keep[63:40] <= 24'h0;
                end else if(stage_join_keep == 40'hffffffffff) begin
                    stage_reinsertion_data[319:0] <= stage_join_data[319:0]; 
                    stage_reinsertion_data[351:320] <= stage_join_crc; 
                    stage_reinsertion_data[511:352] <= 160'b0; 
                    stage_reinsertion_keep[43:0] <= 44'hfffffffffff;
                    stage_reinsertion_keep[63:44] <= 20'h0;
                end else if(stage_join_keep == 44'hfffffffffff) begin 
                    stage_reinsertion_data[351:0] <= stage_join_data[351:0]; 
                    stage_reinsertion_data[383:352] <= stage_join_crc; 
                    stage_reinsertion_data[511:384] <= 128'b0; 
                    stage_reinsertion_keep[47:0] <= 48'hffffffffffff;
                    stage_reinsertion_keep[63:48] <= 16'h0;
                end else if(stage_join_keep == 48'hffffffffffff) begin 
                    stage_reinsertion_data[383:0] <= stage_join_data[383:0]; 
                    stage_reinsertion_data[415:384] <= stage_join_crc; 
                    stage_reinsertion_data[511:416] <= 96'b0; 
                    stage_reinsertion_keep[51:0] <= 52'hfffffffffffff;
                    stage_reinsertion_keep[63:52] <= 12'h0;
                end else if(stage_join_keep == 52'hfffffffffffff) begin
                    stage_reinsertion_data[415:0] <= stage_join_data[415:0]; 
                    stage_reinsertion_data[447:416] <= stage_join_crc; 
                    stage_reinsertion_data[511:448] <= 64'b0; 
                    stage_reinsertion_keep[55:0] <= 56'hffffffffffffff;
                    stage_reinsertion_keep[63:56] <= 8'h0;
                end else if(stage_join_keep == 56'hffffffffffffff) begin
                    stage_reinsertion_data[447:0] <= stage_join_data[447:0]; 
                    stage_reinsertion_data[479:448] <= stage_join_crc; 
                    stage_reinsertion_data[511:480] <= 32'b0; 
                    stage_reinsertion_keep[59:0] <= 60'hfffffffffffffff;
                    stage_reinsertion_keep[63:60] <= 4'h0;
                end else if(stage_join_keep == 60'hfffffffffffffff) begin
                    stage_reinsertion_data[479:0] <= stage_join_data[479:0]; 
                    stage_reinsertion_data[511:480] <= stage_join_crc; 
                    stage_reinsertion_keep[63:0] <= 64'hffffffffffffffff;
                end
            end 

        end


        ///////////////////////////////////////////////////////////////////////
        //
        // STAGE 5: FORMATION OF A NEW WORD (if required)
        //
        ///////////////////////////////////////////////////////////////////////

        // Only act if pipeline is stalled 
        if(stall_pipeline) begin 
            switch_output <= 1; 
            stage_add_word_valid <= 1'b1; 
            stage_add_word_data[31:0] <= stage_reinsertion_crc; 
            stage_add_word_data[511:32] <= 480'b0; 
            stage_add_word_crc <= stage_reinsertion_crc; 
            stage_add_word_keep[3:0] <= 4'hf; 
            stage_add_word_keep[63:4] <= 0; 
            stage_add_word_last <= 1'b1; 
            stall_pipeline <= 1'b0; 
        end else begin 
            switch_output <= 0; 
            stage_add_word_valid <= 1'b0; 
            stage_add_word_data <= 512'b0; 
            stage_add_word_crc <= 32'b0; 
            stage_add_word_keep <= 64'b0; 
            stage_add_word_last <= 1'b1; 
        end 
    end
end 

// Installing an ILA inside the ICRC to check for data
// ila_icrc_pipeline inst_ila_icrc_pipeline(
//     .clk(nclk), 
//     .probe0(stage_masking_valid),           // 1
//     .probe1(d),                             // 512
//     .probe2(pipeline_to_fifo_data),         // 512
//     .probe3(m_axis_rx.tready),              // 1
//     .probe4(m_axis_tx.tready)               // 1
// );


///////////////////////////////////////////////////////////////////////////////////
//
// BUFFER-FIFO AT THE END OF THE PIPELINE
// 
//////////////////////////////////////////////////////////////////////////////////

// Inputs to the FIFO 
assign pipeline_to_fifo_data = switch_output ? stage_add_word_data : stage_reinsertion_data; 
assign pipeline_to_fifo_valid = switch_output ? stage_add_word_valid : stage_reinsertion_valid; 
assign pipeline_to_fifo_last = switch_output ? stage_add_word_last : stage_reinsertion_last; 
assign pipeline_to_fifo_keep = switch_output ? stage_add_word_keep : stage_reinsertion_keep; 
assign pipeline_to_fifo_reset = !nresetn; 


// Initialisation of the FIFO 
buffer_fifo bf(
    .clock(nclk), 
    .reset(pipeline_to_fifo_reset), 
    .input_data(pipeline_to_fifo_data), 
    .input_keep(pipeline_to_fifo_keep), 
    .input_last(pipeline_to_fifo_last), 
    .write_enable(pipeline_to_fifo_valid), 
    .read_enable(m_axis_tx.tready), 
    .output_data(m_axis_tx.tdata), 
    .output_keep(m_axis_tx.tkeep), 
    .output_last(m_axis_tx.tlast), 
    .full(full_signal), 
    .empty(empty_output), 
    .halffull(halffull_signal)
); 

assign m_axis_rx.tready = ~halffull_signal & ~crc32_in_flight_comb & ~full_signal; 
assign m_axis_tx.tvalid = ~empty_output;

/* always_ff @(posedge nclk) begin 
    if(pipeline_to_fifo_reset) begin 
        m_axis_tx.tvalid <= 0; 
    end else begin 
        m_axis_tx.tvalid <= !empty_output; 
    end 
end */ 

//////////////////////////////////////////////////////////////////////////////////
//
// ASSIGN OUTPUTS TO THE PIPELINE
//
//////////////////////////////////////////////////////////////////////////////////

// assign m_axis_tx.tdata = switch_output ? stage_add_word_data : stage_reinsertion_data; 
// assign m_axis_tx.tvalid = switch_output ? stage_add_word_valid : stage_reinsertion_valid; 
// assign m_axis_tx.tlast = switch_output ? stage_add_word_last : stage_reinsertion_last; 
// assign m_axis_tx.tkeep = switch_output ? stage_add_word_keep : stage_reinsertion_keep; 


////////////////////////////////////////////////////////////////////////////////////
//
// ASSIGN READY INPUT TO THE PIPELINE
//
////////////////////////////////////////////////////////////////////////////////////

// assign m_axis_rx.tready = m_axis_tx.tready; 

endmodule