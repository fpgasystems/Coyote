
`timescale 1ns / 1ps

import lynxTypes::*;

/**
 * @brief  HBM AXI split
 *
 * Splits 512-bit AXI sink to 2x 256-bit AXI sources
 */
/*
module hbm_split (
    input  logic                aclk,
    input  logic                aresetn,

    AXI4.s                      axi_in,
    AXI4.m                      axi_out [2]
);

AXI4 #(.AXI4_DATA_BITS)
    
endmodule*/