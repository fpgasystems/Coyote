

// this is a simple pass through
arrow_top arrow_top_inst(
    // AXI4L CONTROL
    .axi_ctrl(axi_ctrl),

    // NOTIFY
    .notify(notify),

    // DESCRIPTORS
    .sq_rd(sq_rd),
    .sq_wr(sq_wr),
    .cq_rd(cq_rd),
    .cq_wr(cq_wr),
    .rq_rd(rq_rd),
    .rq_wr(rq_wr),

    // HOST DATA STREAMS
    .axis_host_recv(axis_host_recv),
    .axis_host_send(axis_host_send),

    // RDMA DATA STREAMS REQUESTER
    .axis_rreq_recv(axis_rreq_recv),
    .axis_rreq_send(axis_rreq_send),

    // RDMA DATA STREAMS RESPONDER
    .axis_rrsp_recv(axis_rrsp_recv),
    .axis_rrsp_send(axis_rrsp_send),

    // Clock and reset
    .aclk(aclk),
    .aresetn(aresetn)
);//*/

`ifndef XILINX_SIMULATOR
    ila_ctrl inst_ila_ctrl (
        .probe0(axi_ctrl.araddr),
        .probe1(axi_ctrl.arprot),
        .probe2(axi_ctrl.arqos),
        .probe3(axi_ctrl.arregion),
        .probe4(axi_ctrl.arready),
        .probe5(axi_ctrl.arvalid),
        .probe6(axi_ctrl.awaddr),
        .probe7(axi_ctrl.awprot),
        .probe8(axi_ctrl.awqos),
        .probe9(axi_ctrl.awregion),
        .probe10(axi_ctrl.awready),
        .probe11(axi_ctrl.awvalid),
        .probe12(axi_ctrl.rdata),
        .probe13(axi_ctrl.rresp),
        .probe14(axi_ctrl.rready),
        .probe15(axi_ctrl.rvalid),
        .probe16(axi_ctrl.wdata),
        .probe17(axi_ctrl.wstrb),
        .probe18(axi_ctrl.wready),
        .probe19(axi_ctrl.wvalid),
        .probe20(axi_ctrl.bresp),
        .probe21(axi_ctrl.bready),
        .probe22(axi_ctrl.bvalid),
        .probe23(notify.data.pid),
        .probe24(notify.data.value),
        .probe25(notify.valid),
        .probe26(notify.ready),
        .probe27(sq_rd.data.opcode),
        .probe28(sq_rd.data.strm),
        .probe29(sq_rd.data.mode),
        .probe30(sq_rd.data.rdma),
        .probe31(sq_rd.data.remote),
        .probe32(sq_rd.data.vfid),
        .probe33(sq_rd.data.pid),
        .probe34(sq_rd.data.dest),
        .probe35(sq_rd.data.last),
        .probe36(sq_rd.data.vaddr),
        .probe37(sq_rd.data.len),
        .probe38(sq_rd.data.actv),
        .probe39(sq_rd.data.host),
        .probe40(sq_rd.data.offs),
        .probe41(sq_rd.valid),
        .probe42(sq_rd.ready),
        .probe43(sq_wr.data.opcode),
        .probe44(sq_wr.data.strm),
        .probe45(sq_wr.data.mode),
        .probe46(sq_wr.data.rdma),
        .probe47(sq_wr.data.remote),
        .probe48(sq_wr.data.vfid),
        .probe49(sq_wr.data.pid),
        .probe50(sq_wr.data.dest),
        .probe51(sq_wr.data.last),
        .probe52(sq_wr.data.vaddr),
        .probe53(sq_wr.data.len),
        .probe54(sq_wr.data.actv),
        .probe55(sq_wr.data.host),
        .probe56(sq_wr.data.offs),
        .probe57(sq_wr.valid),
        .probe58(sq_wr.ready),
        .probe59(cq_rd.data.opcode),
        .probe60(cq_rd.data.strm),
        .probe61(cq_rd.data.remote),
        .probe62(cq_rd.data.host),
        .probe63(cq_rd.data.dest),
        .probe64(cq_rd.data.pid),
        .probe65(cq_rd.data.vfid),
        .probe66(cq_rd.valid),
        .probe67(cq_rd.ready),
        .probe68(cq_wr.data.opcode),
        .probe69(cq_wr.data.strm),
        .probe70(cq_wr.data.remote),
        .probe71(cq_wr.data.host),
        .probe72(cq_wr.data.dest),
        .probe73(cq_wr.data.pid),
        .probe74(cq_wr.data.vfid),
        .probe75(cq_wr.valid),
        .probe76(cq_wr.ready),
        .probe77(rq_wr.data.opcode),
        .probe78(rq_wr.data.strm),
        .probe79(rq_wr.data.mode),
        .probe80(rq_wr.data.rdma),
        .probe81(rq_wr.data.remote),
        .probe82(rq_wr.data.vfid),
        .probe83(rq_wr.data.pid),
        .probe84(rq_wr.data.dest),
        .probe85(rq_wr.data.last),
        .probe86(rq_wr.data.vaddr),
        .probe87(rq_wr.data.len),
        .probe88(rq_wr.data.actv),
        .probe89(rq_wr.data.host),
        .probe90(rq_wr.data.offs),
        .probe91(rq_wr.valid),
        .probe92(rq_wr.ready),
        .probe93(rq_rd.data.opcode),
        .probe94(rq_rd.data.strm),
        .probe95(rq_rd.data.mode),
        .probe96(rq_rd.data.rdma),
        .probe97(rq_rd.data.remote),
        .probe98(rq_rd.data.vfid),
        .probe99(rq_rd.data.pid),
        .probe100(rq_rd.data.dest),
        .probe101(rq_rd.data.last),
        .probe102(rq_rd.data.vaddr),
        .probe103(rq_rd.data.len),
        .probe104(rq_rd.data.actv),
        .probe105(rq_rd.data.host),
        .probe106(rq_rd.data.offs),
        .probe107(rq_rd.valid),
        .probe108(rq_rd.ready),
        .probe109(axis_host_recv[0].tdata),
        .probe110(axis_host_recv[0].tkeep),
        .probe111(axis_host_recv[0].tlast),
        .probe112(axis_host_recv[0].tready),
        .probe113(axis_host_recv[0].tvalid),
        .probe114(axis_host_recv[1].tdata),
        .probe115(axis_host_recv[1].tkeep),
        .probe116(axis_host_recv[1].tlast),
        .probe117(axis_host_recv[1].tready),
        .probe118(axis_host_recv[1].tvalid),
        .probe119(axis_host_send[0].tdata),
        .probe120(axis_host_send[0].tkeep),
        .probe121(axis_host_send[0].tlast),
        .probe122(axis_host_send[0].tready),
        .probe123(axis_host_send[0].tvalid),
        .probe124(axis_host_send[1].tdata),
        .probe125(axis_host_send[1].tkeep),
        .probe126(axis_host_send[1].tlast),
        .probe127(axis_host_send[1].tready),
        .probe128(axis_host_send[1].tvalid),
        .probe129(axis_rreq_recv[0].tdata),
        .probe130(axis_rreq_recv[0].tkeep),
        .probe131(axis_rreq_recv[0].tlast),
        .probe132(axis_rreq_recv[0].tready),
        .probe133(axis_rreq_recv[0].tvalid),
        .probe134(axis_rreq_send[0].tdata),
        .probe135(axis_rreq_send[0].tkeep),
        .probe136(axis_rreq_send[0].tlast),
        .probe137(axis_rreq_send[0].tready),
        .probe138(axis_rreq_send[0].tvalid),
        .probe139(axis_rrsp_recv[0].tdata),
        .probe140(axis_rrsp_recv[0].tkeep),
        .probe141(axis_rrsp_recv[0].tlast),
        .probe142(axis_rrsp_recv[0].tready),
        .probe143(axis_rrsp_recv[0].tvalid),
        .probe144(axis_rrsp_send[0].tdata),
        .probe145(axis_rrsp_send[0].tkeep),
        .probe146(axis_rrsp_send[0].tlast),
        .probe147(axis_rrsp_send[0].tready),
        .probe148(axis_rrsp_send[0].tvalid),
        .clk(aclk)
    );

`endif
