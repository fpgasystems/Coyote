-------------------------------------------------------------------------------
-- MSB-first 64b CRC32, generator 0x1EDC6F41
--
-- Copyright (c) 2022 ETH Zurich.
-- All rights reserved.
--
-- This file is distributed under the terms in the attached LICENSE file.
-- If you do not find this file, copies can be found by writing to:
-- ETH Zurich D-INFK, Stampfenbachstrasse 114, CH-8092 Zurich. Attn: Systems Group
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity crc_64_32_1edc6f41 is
port (
    R   :  in std_logic_vector(31 downto 0);
    X   :  in std_logic_vector(63 downto 0);
    R_n : out std_logic_vector(31 downto 0)
);
end crc_64_32_1edc6f41;

architecture functional of crc_64_32_1edc6f41 is
begin

R_n(31) <= X(3) xor X(4) xor X(5) xor X(6) xor X(7) xor X(8) xor X(11) xor X(15) xor X(16) xor X(17) xor X(20) xor X(22) xor X(24) xor X(25) xor X(26) xor X(27) xor X(29) xor X(30) xor X(34) xor X(35) xor X(36) xor X(41) xor X(42) xor X(44) xor X(45) xor X(46) xor X(47) xor X(50) xor X(52) xor X(53) xor X(58) xor X(61) xor X(63) xor R(2) xor R(3) xor R(4) xor R(9) xor R(10) xor R(12) xor R(13) xor R(14) xor R(15) xor R(18) xor R(20) xor R(21) xor R(26) xor R(29) xor R(31) ;
R_n(30) <= X(2) xor X(3) xor X(4) xor X(5) xor X(6) xor X(7) xor X(10) xor X(14) xor X(15) xor X(16) xor X(19) xor X(21) xor X(23) xor X(24) xor X(25) xor X(26) xor X(28) xor X(29) xor X(33) xor X(34) xor X(35) xor X(40) xor X(41) xor X(43) xor X(44) xor X(45) xor X(46) xor X(49) xor X(51) xor X(52) xor X(57) xor X(60) xor X(62) xor X(63) xor R(1) xor R(2) xor R(3) xor R(8) xor R(9) xor R(11) xor R(12) xor R(13) xor R(14) xor R(17) xor R(19) xor R(20) xor R(25) xor R(28) xor R(30) xor R(31) ;
R_n(29) <= X(1) xor X(2) xor X(3) xor X(4) xor X(5) xor X(6) xor X(9) xor X(13) xor X(14) xor X(15) xor X(18) xor X(20) xor X(22) xor X(23) xor X(24) xor X(25) xor X(27) xor X(28) xor X(32) xor X(33) xor X(34) xor X(39) xor X(40) xor X(42) xor X(43) xor X(44) xor X(45) xor X(48) xor X(50) xor X(51) xor X(56) xor X(59) xor X(61) xor X(62) xor X(63) xor R(0) xor R(1) xor R(2) xor R(7) xor R(8) xor R(10) xor R(11) xor R(12) xor R(13) xor R(16) xor R(18) xor R(19) xor R(24) xor R(27) xor R(29) xor R(30) xor R(31) ;
R_n(28) <= X(0) xor X(1) xor X(2) xor X(3) xor X(4) xor X(5) xor X(8) xor X(12) xor X(13) xor X(14) xor X(17) xor X(19) xor X(21) xor X(22) xor X(23) xor X(24) xor X(26) xor X(27) xor X(31) xor X(32) xor X(33) xor X(38) xor X(39) xor X(41) xor X(42) xor X(43) xor X(44) xor X(47) xor X(49) xor X(50) xor X(55) xor X(58) xor X(60) xor X(61) xor X(62) xor R(0) xor R(1) xor R(6) xor R(7) xor R(9) xor R(10) xor R(11) xor R(12) xor R(15) xor R(17) xor R(18) xor R(23) xor R(26) xor R(28) xor R(29) xor R(30) ;
R_n(27) <= X(0) xor X(1) xor X(2) xor X(5) xor X(6) xor X(8) xor X(12) xor X(13) xor X(15) xor X(17) xor X(18) xor X(21) xor X(23) xor X(24) xor X(27) xor X(29) xor X(31) xor X(32) xor X(34) xor X(35) xor X(36) xor X(37) xor X(38) xor X(40) xor X(43) xor X(44) xor X(45) xor X(47) xor X(48) xor X(49) xor X(50) xor X(52) xor X(53) xor X(54) xor X(57) xor X(58) xor X(59) xor X(60) xor R(0) xor R(2) xor R(3) xor R(4) xor R(5) xor R(6) xor R(8) xor R(11) xor R(12) xor R(13) xor R(15) xor R(16) xor R(17) xor R(18) xor R(20) xor R(21) xor R(22) xor R(25) xor R(26) xor R(27) xor R(28) ;
R_n(26) <= X(0) xor X(1) xor X(3) xor X(6) xor X(8) xor X(12) xor X(14) xor X(15) xor X(23) xor X(24) xor X(25) xor X(27) xor X(28) xor X(29) xor X(31) xor X(33) xor X(37) xor X(39) xor X(41) xor X(43) xor X(45) xor X(48) xor X(49) xor X(50) xor X(51) xor X(56) xor X(57) xor X(59) xor X(61) xor X(63) xor R(1) xor R(5) xor R(7) xor R(9) xor R(11) xor R(13) xor R(16) xor R(17) xor R(18) xor R(19) xor R(24) xor R(25) xor R(27) xor R(29) xor R(31) ;
R_n(25) <= X(0) xor X(2) xor X(3) xor X(4) xor X(6) xor X(8) xor X(13) xor X(14) xor X(15) xor X(16) xor X(17) xor X(20) xor X(23) xor X(25) xor X(28) xor X(29) xor X(32) xor X(34) xor X(35) xor X(38) xor X(40) xor X(41) xor X(45) xor X(46) xor X(48) xor X(49) xor X(52) xor X(53) xor X(55) xor X(56) xor X(60) xor X(61) xor X(62) xor R(0) xor R(2) xor R(3) xor R(6) xor R(8) xor R(9) xor R(13) xor R(14) xor R(16) xor R(17) xor R(20) xor R(21) xor R(23) xor R(24) xor R(28) xor R(29) xor R(30) ;
R_n(24) <= X(1) xor X(2) xor X(4) xor X(6) xor X(8) xor X(11) xor X(12) xor X(13) xor X(14) xor X(17) xor X(19) xor X(20) xor X(25) xor X(26) xor X(28) xor X(29) xor X(30) xor X(31) xor X(33) xor X(35) xor X(36) xor X(37) xor X(39) xor X(40) xor X(41) xor X(42) xor X(46) xor X(48) xor X(50) xor X(51) xor X(53) xor X(54) xor X(55) xor X(58) xor X(59) xor X(60) xor R(1) xor R(3) xor R(4) xor R(5) xor R(7) xor R(8) xor R(9) xor R(10) xor R(14) xor R(16) xor R(18) xor R(19) xor R(21) xor R(22) xor R(23) xor R(26) xor R(27) xor R(28) ;
R_n(23) <= X(0) xor X(1) xor X(3) xor X(5) xor X(7) xor X(10) xor X(11) xor X(12) xor X(13) xor X(16) xor X(18) xor X(19) xor X(24) xor X(25) xor X(27) xor X(28) xor X(29) xor X(30) xor X(32) xor X(34) xor X(35) xor X(36) xor X(38) xor X(39) xor X(40) xor X(41) xor X(45) xor X(47) xor X(49) xor X(50) xor X(52) xor X(53) xor X(54) xor X(57) xor X(58) xor X(59) xor X(63) xor R(0) xor R(2) xor R(3) xor R(4) xor R(6) xor R(7) xor R(8) xor R(9) xor R(13) xor R(15) xor R(17) xor R(18) xor R(20) xor R(21) xor R(22) xor R(25) xor R(26) xor R(27) xor R(31) ;
R_n(22) <= X(0) xor X(2) xor X(3) xor X(5) xor X(7) xor X(8) xor X(9) xor X(10) xor X(12) xor X(16) xor X(18) xor X(20) xor X(22) xor X(23) xor X(25) xor X(28) xor X(30) xor X(31) xor X(33) xor X(36) xor X(37) xor X(38) xor X(39) xor X(40) xor X(41) xor X(42) xor X(45) xor X(47) xor X(48) xor X(49) xor X(50) xor X(51) xor X(56) xor X(57) xor X(61) xor X(62) xor R(1) xor R(4) xor R(5) xor R(6) xor R(7) xor R(8) xor R(9) xor R(10) xor R(13) xor R(15) xor R(16) xor R(17) xor R(18) xor R(19) xor R(24) xor R(25) xor R(29) xor R(30) ;
R_n(21) <= X(1) xor X(2) xor X(3) xor X(5) xor X(9) xor X(16) xor X(19) xor X(20) xor X(21) xor X(25) xor X(26) xor X(32) xor X(34) xor X(37) xor X(38) xor X(39) xor X(40) xor X(42) xor X(45) xor X(48) xor X(49) xor X(52) xor X(53) xor X(55) xor X(56) xor X(58) xor X(60) xor X(63) xor R(0) xor R(2) xor R(5) xor R(6) xor R(7) xor R(8) xor R(10) xor R(13) xor R(16) xor R(17) xor R(20) xor R(21) xor R(23) xor R(24) xor R(26) xor R(28) xor R(31) ;
R_n(20) <= X(0) xor X(1) xor X(2) xor X(4) xor X(8) xor X(15) xor X(18) xor X(19) xor X(20) xor X(24) xor X(25) xor X(31) xor X(33) xor X(36) xor X(37) xor X(38) xor X(39) xor X(41) xor X(44) xor X(47) xor X(48) xor X(51) xor X(52) xor X(54) xor X(55) xor X(57) xor X(59) xor X(62) xor X(63) xor R(1) xor R(4) xor R(5) xor R(6) xor R(7) xor R(9) xor R(12) xor R(15) xor R(16) xor R(19) xor R(20) xor R(22) xor R(23) xor R(25) xor R(27) xor R(30) xor R(31) ;
R_n(19) <= X(0) xor X(1) xor X(4) xor X(5) xor X(6) xor X(8) xor X(11) xor X(14) xor X(15) xor X(16) xor X(18) xor X(19) xor X(20) xor X(22) xor X(23) xor X(25) xor X(26) xor X(27) xor X(29) xor X(32) xor X(34) xor X(37) xor X(38) xor X(40) xor X(41) xor X(42) xor X(43) xor X(44) xor X(45) xor X(51) xor X(52) xor X(54) xor X(56) xor X(62) xor X(63) xor R(0) xor R(2) xor R(5) xor R(6) xor R(8) xor R(9) xor R(10) xor R(11) xor R(12) xor R(13) xor R(19) xor R(20) xor R(22) xor R(24) xor R(30) xor R(31) ;
R_n(18) <= X(0) xor X(6) xor X(8) xor X(10) xor X(11) xor X(13) xor X(14) xor X(16) xor X(18) xor X(19) xor X(20) xor X(21) xor X(27) xor X(28) xor X(29) xor X(30) xor X(31) xor X(33) xor X(34) xor X(35) xor X(37) xor X(39) xor X(40) xor X(43) xor X(45) xor X(46) xor X(47) xor X(51) xor X(52) xor X(55) xor X(58) xor X(62) xor X(63) xor R(1) xor R(2) xor R(3) xor R(5) xor R(7) xor R(8) xor R(11) xor R(13) xor R(14) xor R(15) xor R(19) xor R(20) xor R(23) xor R(26) xor R(30) xor R(31) ;
R_n(17) <= X(3) xor X(4) xor X(6) xor X(8) xor X(9) xor X(10) xor X(11) xor X(12) xor X(13) xor X(16) xor X(18) xor X(19) xor X(22) xor X(24) xor X(25) xor X(28) xor X(32) xor X(33) xor X(35) xor X(38) xor X(39) xor X(41) xor X(47) xor X(51) xor X(52) xor X(53) xor X(54) xor X(57) xor X(58) xor X(62) xor X(63) xor R(0) xor R(1) xor R(3) xor R(6) xor R(7) xor R(9) xor R(15) xor R(19) xor R(20) xor R(21) xor R(22) xor R(25) xor R(26) xor R(30) xor R(31) ;
R_n(16) <= X(2) xor X(3) xor X(5) xor X(7) xor X(8) xor X(9) xor X(10) xor X(11) xor X(12) xor X(15) xor X(17) xor X(18) xor X(21) xor X(23) xor X(24) xor X(27) xor X(31) xor X(32) xor X(34) xor X(37) xor X(38) xor X(40) xor X(46) xor X(50) xor X(51) xor X(52) xor X(53) xor X(56) xor X(57) xor X(61) xor X(62) xor R(0) xor R(2) xor R(5) xor R(6) xor R(8) xor R(14) xor R(18) xor R(19) xor R(20) xor R(21) xor R(24) xor R(25) xor R(29) xor R(30) ;
R_n(15) <= X(1) xor X(2) xor X(4) xor X(6) xor X(7) xor X(8) xor X(9) xor X(10) xor X(11) xor X(14) xor X(16) xor X(17) xor X(20) xor X(22) xor X(23) xor X(26) xor X(30) xor X(31) xor X(33) xor X(36) xor X(37) xor X(39) xor X(45) xor X(49) xor X(50) xor X(51) xor X(52) xor X(55) xor X(56) xor X(60) xor X(61) xor R(1) xor R(4) xor R(5) xor R(7) xor R(13) xor R(17) xor R(18) xor R(19) xor R(20) xor R(23) xor R(24) xor R(28) xor R(29) ;
R_n(14) <= X(0) xor X(1) xor X(3) xor X(5) xor X(6) xor X(7) xor X(8) xor X(9) xor X(10) xor X(13) xor X(15) xor X(16) xor X(19) xor X(21) xor X(22) xor X(25) xor X(29) xor X(30) xor X(32) xor X(35) xor X(36) xor X(38) xor X(44) xor X(48) xor X(49) xor X(50) xor X(51) xor X(54) xor X(55) xor X(59) xor X(60) xor R(0) xor R(3) xor R(4) xor R(6) xor R(12) xor R(16) xor R(17) xor R(18) xor R(19) xor R(22) xor R(23) xor R(27) xor R(28) ;
R_n(13) <= X(0) xor X(2) xor X(3) xor X(9) xor X(11) xor X(12) xor X(14) xor X(16) xor X(17) xor X(18) xor X(21) xor X(22) xor X(25) xor X(26) xor X(27) xor X(28) xor X(30) xor X(31) xor X(36) xor X(37) xor X(41) xor X(42) xor X(43) xor X(44) xor X(45) xor X(46) xor X(48) xor X(49) xor X(52) xor X(54) xor X(59) xor X(61) xor X(63) xor R(4) xor R(5) xor R(9) xor R(10) xor R(11) xor R(12) xor R(13) xor R(14) xor R(16) xor R(17) xor R(20) xor R(22) xor R(27) xor R(29) xor R(31) ;
R_n(12) <= X(1) xor X(2) xor X(3) xor X(4) xor X(5) xor X(6) xor X(7) xor X(10) xor X(13) xor X(21) xor X(22) xor X(34) xor X(40) xor X(43) xor X(46) xor X(48) xor X(50) xor X(51) xor X(52) xor X(60) xor X(61) xor X(62) xor X(63) xor R(2) xor R(8) xor R(11) xor R(14) xor R(16) xor R(18) xor R(19) xor R(20) xor R(28) xor R(29) xor R(30) xor R(31) ;
R_n(11) <= X(0) xor X(1) xor X(2) xor X(3) xor X(4) xor X(5) xor X(6) xor X(9) xor X(12) xor X(20) xor X(21) xor X(33) xor X(39) xor X(42) xor X(45) xor X(47) xor X(49) xor X(50) xor X(51) xor X(59) xor X(60) xor X(61) xor X(62) xor X(63) xor R(1) xor R(7) xor R(10) xor R(13) xor R(15) xor R(17) xor R(18) xor R(19) xor R(27) xor R(28) xor R(29) xor R(30) xor R(31) ;
R_n(10) <= X(0) xor X(1) xor X(2) xor X(6) xor X(7) xor X(15) xor X(16) xor X(17) xor X(19) xor X(22) xor X(24) xor X(25) xor X(26) xor X(27) xor X(29) xor X(30) xor X(32) xor X(34) xor X(35) xor X(36) xor X(38) xor X(42) xor X(45) xor X(47) xor X(48) xor X(49) xor X(52) xor X(53) xor X(59) xor X(60) xor X(62) xor X(63) xor R(0) xor R(2) xor R(3) xor R(4) xor R(6) xor R(10) xor R(13) xor R(15) xor R(16) xor R(17) xor R(20) xor R(21) xor R(27) xor R(28) xor R(30) xor R(31) ;
R_n(9) <= X(0) xor X(1) xor X(3) xor X(4) xor X(7) xor X(8) xor X(11) xor X(14) xor X(17) xor X(18) xor X(20) xor X(21) xor X(22) xor X(23) xor X(27) xor X(28) xor X(30) xor X(31) xor X(33) xor X(36) xor X(37) xor X(42) xor X(45) xor X(48) xor X(50) xor X(51) xor X(53) xor X(59) xor X(62) xor R(1) xor R(4) xor R(5) xor R(10) xor R(13) xor R(16) xor R(18) xor R(19) xor R(21) xor R(27) xor R(30) ;
R_n(8) <= X(0) xor X(2) xor X(4) xor X(5) xor X(8) xor X(10) xor X(11) xor X(13) xor X(15) xor X(19) xor X(21) xor X(24) xor X(25) xor X(32) xor X(34) xor X(42) xor X(45) xor X(46) xor X(49) xor X(53) xor R(0) xor R(2) xor R(10) xor R(13) xor R(14) xor R(17) xor R(21) ;
R_n(7) <= X(1) xor X(5) xor X(6) xor X(8) xor X(9) xor X(10) xor X(11) xor X(12) xor X(14) xor X(15) xor X(16) xor X(17) xor X(18) xor X(22) xor X(23) xor X(25) xor X(26) xor X(27) xor X(29) xor X(30) xor X(31) xor X(33) xor X(34) xor X(35) xor X(36) xor X(42) xor X(46) xor X(47) xor X(48) xor X(50) xor X(53) xor X(58) xor X(61) xor X(63) xor R(1) xor R(2) xor R(3) xor R(4) xor R(10) xor R(14) xor R(15) xor R(16) xor R(18) xor R(21) xor R(26) xor R(29) xor R(31) ;
R_n(6) <= X(0) xor X(4) xor X(5) xor X(7) xor X(8) xor X(9) xor X(10) xor X(11) xor X(13) xor X(14) xor X(15) xor X(16) xor X(17) xor X(21) xor X(22) xor X(24) xor X(25) xor X(26) xor X(28) xor X(29) xor X(30) xor X(32) xor X(33) xor X(34) xor X(35) xor X(41) xor X(45) xor X(46) xor X(47) xor X(49) xor X(52) xor X(57) xor X(60) xor X(62) xor R(0) xor R(1) xor R(2) xor R(3) xor R(9) xor R(13) xor R(14) xor R(15) xor R(17) xor R(20) xor R(25) xor R(28) xor R(30) ;
R_n(5) <= X(5) xor X(9) xor X(10) xor X(11) xor X(12) xor X(13) xor X(14) xor X(17) xor X(21) xor X(22) xor X(23) xor X(26) xor X(28) xor X(30) xor X(31) xor X(32) xor X(33) xor X(35) xor X(36) xor X(40) xor X(41) xor X(42) xor X(47) xor X(48) xor X(50) xor X(51) xor X(52) xor X(53) xor X(56) xor X(58) xor X(59) xor R(0) xor R(1) xor R(3) xor R(4) xor R(8) xor R(9) xor R(10) xor R(15) xor R(16) xor R(18) xor R(19) xor R(20) xor R(21) xor R(24) xor R(26) xor R(27) ;
R_n(4) <= X(4) xor X(8) xor X(9) xor X(10) xor X(11) xor X(12) xor X(13) xor X(16) xor X(20) xor X(21) xor X(22) xor X(25) xor X(27) xor X(29) xor X(30) xor X(31) xor X(32) xor X(34) xor X(35) xor X(39) xor X(40) xor X(41) xor X(46) xor X(47) xor X(49) xor X(50) xor X(51) xor X(52) xor X(55) xor X(57) xor X(58) xor X(63) xor R(0) xor R(2) xor R(3) xor R(7) xor R(8) xor R(9) xor R(14) xor R(15) xor R(17) xor R(18) xor R(19) xor R(20) xor R(23) xor R(25) xor R(26) xor R(31) ;
R_n(3) <= X(3) xor X(7) xor X(8) xor X(9) xor X(10) xor X(11) xor X(12) xor X(15) xor X(19) xor X(20) xor X(21) xor X(24) xor X(26) xor X(28) xor X(29) xor X(30) xor X(31) xor X(33) xor X(34) xor X(38) xor X(39) xor X(40) xor X(45) xor X(46) xor X(48) xor X(49) xor X(50) xor X(51) xor X(54) xor X(56) xor X(57) xor X(62) xor R(1) xor R(2) xor R(6) xor R(7) xor R(8) xor R(13) xor R(14) xor R(16) xor R(17) xor R(18) xor R(19) xor R(22) xor R(24) xor R(25) xor R(30) ;
R_n(2) <= X(2) xor X(6) xor X(7) xor X(8) xor X(9) xor X(10) xor X(11) xor X(14) xor X(18) xor X(19) xor X(20) xor X(23) xor X(25) xor X(27) xor X(28) xor X(29) xor X(30) xor X(32) xor X(33) xor X(37) xor X(38) xor X(39) xor X(44) xor X(45) xor X(47) xor X(48) xor X(49) xor X(50) xor X(53) xor X(55) xor X(56) xor X(61) xor R(0) xor R(1) xor R(5) xor R(6) xor R(7) xor R(12) xor R(13) xor R(15) xor R(16) xor R(17) xor R(18) xor R(21) xor R(23) xor R(24) xor R(29) ;
R_n(1) <= X(1) xor X(5) xor X(6) xor X(7) xor X(8) xor X(9) xor X(10) xor X(13) xor X(17) xor X(18) xor X(19) xor X(22) xor X(24) xor X(26) xor X(27) xor X(28) xor X(29) xor X(31) xor X(32) xor X(36) xor X(37) xor X(38) xor X(43) xor X(44) xor X(46) xor X(47) xor X(48) xor X(49) xor X(52) xor X(54) xor X(55) xor X(60) xor X(63) xor R(0) xor R(4) xor R(5) xor R(6) xor R(11) xor R(12) xor R(14) xor R(15) xor R(16) xor R(17) xor R(20) xor R(22) xor R(23) xor R(28) xor R(31) ;
R_n(0) <= X(0) xor X(4) xor X(5) xor X(6) xor X(7) xor X(8) xor X(9) xor X(12) xor X(16) xor X(17) xor X(18) xor X(21) xor X(23) xor X(25) xor X(26) xor X(27) xor X(28) xor X(30) xor X(31) xor X(35) xor X(36) xor X(37) xor X(42) xor X(43) xor X(45) xor X(46) xor X(47) xor X(48) xor X(51) xor X(53) xor X(54) xor X(59) xor X(62) xor R(3) xor R(4) xor R(5) xor R(10) xor R(11) xor R(13) xor R(14) xor R(15) xor R(16) xor R(19) xor R(21) xor R(22) xor R(27) xor R(30) ;

end functional;
