localparam [7:0]
	OPCODE_SETUPPEER  = 17,
	OPCODE_ADDPEER    = 18,
	OPCODE_REMOVEPEER = 19,
	OPCODE_SETLEADER  = 20,

	OPCODE_SETCOMMITCNT  = 25,
	OPCODE_SETSILENCECNT = 26,
	OPCODE_SETHTSIZE     = 27,

	OPCODE_TOGGLEDEAD = 28,

	OPCODE_SYNCDRAM = 29,

	OPCODE_READREQ    = 0,
	OPCODE_WRITEREQ   = 1,
	OPCODE_PROPOSAL   = 2,
	OPCODE_ACKPROPOSE = 3,
	OPCODE_COMMIT     = 4,
	OPCODE_SYNCREQ    = 5,
	OPCODE_SYNCRESP   = 6,
	OPCODE_SYNCCOMMIT = 7,

	OPCODE_UNVERSIONEDWRITE = 31,		
	OPCODE_UNVERSIONEDDELETE = 47,

	OPCODE_READCONDITIONAL = 64,

    OPCODE_FLUSHDATASTORE = 255,

	OPCODE_DELWRITEREQ   = 32 + 1,
	OPCODE_DELPROPOSAL   = 32 + 2,
	OPCODE_DELACKPROPOSE = 32 + 3,

	OPCODE_CUREPOCH   = 8,
	OPCODE_NEWEPOCH   = 9,
	OPCODE_ACKEPOCH   = 10,
	OPCODE_SYNCLEADER = 11;

localparam [3:0] 
	HTOP_IGNORE = 0,
	HTOP_GET = 1,
	HTOP_SETNEXT = 2,
	HTOP_DELCUR = 3,	
	HTOP_FLIPPOINT = 4,
	HTOP_SETCUR = 5,
	HTOP_GETRAW = 6,
	HTOP_IGNOREPROP = 7,
	HTOP_GETCOND = 8,
	HTOP_FLUSH = 4'hF, //(truncated from 8'hFF)

	HTOP_PRE_INCR = 13, //DEDUP ONLY
	HTOP_PRE_DECR = 14, //DEDUP ONLY


	// these are not supported:
	HTOP_SCAN = 9,
	HTOP_SCANCOND = 10;