
test_top test_top_inst (
    .axi_ctrl(axi_ctrl),
    .notify(notify),
    .sq_rd(sq_rd),
    .sq_wr(sq_wr),
    .cq_rd(cq_rd),
    .cq_wr(cq_wr),
    .axis_host_recv(axis_host_recv),
    .axis_host_send(axis_host_send),
    .aclk(aclk),
    .aresetn(aresetn)
);

`ifndef XILINX_SIMULATOR
ila_ctrl inst_ila_ctrl (
    .probe0(axi_ctrl.araddr),
    .probe1(axi_ctrl.arprot),
    .probe2(axi_ctrl.arqos),
    .probe3(axi_ctrl.arregion),
    .probe4(axi_ctrl.arready),
    .probe5(axi_ctrl.arvalid),
    .probe6(axi_ctrl.awaddr),
    .probe7(axi_ctrl.awprot),
    .probe8(axi_ctrl.awqos),
    .probe9(axi_ctrl.awregion),
    .probe10(axi_ctrl.awready),
    .probe11(axi_ctrl.awvalid),
    .probe12(axi_ctrl.rdata),
    .probe13(axi_ctrl.rresp),
    .probe14(axi_ctrl.rready),
    .probe15(axi_ctrl.rvalid),
    .probe16(axi_ctrl.wdata),
    .probe17(axi_ctrl.wstrb),
    .probe18(axi_ctrl.wready),
    .probe19(axi_ctrl.wvalid),
    .probe20(axi_ctrl.bresp),
    .probe21(axi_ctrl.bready),
    .probe22(axi_ctrl.bvalid),
    .probe23(sq_rd.data.opcode),
    .probe24(sq_rd.data.strm),
    .probe25(sq_rd.data.mode),
    .probe26(sq_rd.data.rdma),
    .probe27(sq_rd.data.remote),
    .probe28(sq_rd.data.vfid),
    .probe29(sq_rd.data.pid),
    .probe30(sq_rd.data.dest),
    .probe31(sq_rd.data.last),
    .probe32(sq_rd.data.vaddr),
    .probe33(sq_rd.data.len),
    .probe34(sq_rd.data.actv),
    .probe35(sq_rd.data.host),
    .probe36(sq_rd.data.offs),
    .probe37(sq_rd.valid),
    .probe38(sq_rd.ready),
    .probe39(sq_wr.data.opcode),
    .probe40(sq_wr.data.strm),
    .probe41(sq_wr.data.mode),
    .probe42(sq_wr.data.rdma),
    .probe43(sq_wr.data.remote),
    .probe44(sq_wr.data.vfid),
    .probe45(sq_wr.data.pid),
    .probe46(sq_wr.data.dest),
    .probe47(sq_wr.data.last),
    .probe48(sq_wr.data.vaddr),
    .probe49(sq_wr.data.len),
    .probe50(sq_wr.data.actv),
    .probe51(sq_wr.data.host),
    .probe52(sq_wr.data.offs),
    .probe53(sq_wr.valid),
    .probe54(sq_wr.ready),
    .probe55(cq_rd.data.opcode),
    .probe56(cq_rd.data.strm),
    .probe57(cq_rd.data.remote),
    .probe58(cq_rd.data.host),
    .probe59(cq_rd.data.dest),
    .probe60(cq_rd.data.pid),
    .probe61(cq_rd.data.vfid),
    .probe62(cq_rd.valid),
    .probe63(cq_rd.ready),
    .probe64(cq_wr.data.opcode),
    .probe65(cq_wr.data.strm),
    .probe66(cq_wr.data.remote),
    .probe67(cq_wr.data.host),
    .probe68(cq_wr.data.dest),
    .probe69(cq_wr.data.pid),
    .probe70(cq_wr.data.vfid),
    .probe71(cq_wr.valid),
    .probe72(cq_wr.ready),
    .probe73(axis_host_recv[0].tdata),
    .probe74(axis_host_recv[0].tkeep),
    .probe75(axis_host_recv[0].tlast),
    .probe76(axis_host_recv[0].tready),
    .probe77(axis_host_recv[0].tvalid),
    .probe78(axis_host_recv[1].tdata),
    .probe79(axis_host_recv[1].tkeep),
    .probe80(axis_host_recv[1].tlast),
    .probe81(axis_host_recv[1].tready),
    .probe82(axis_host_recv[1].tvalid),
    .probe83(axis_host_send[0].tdata),
    .probe84(axis_host_send[0].tkeep),
    .probe85(axis_host_send[0].tlast),
    .probe86(axis_host_send[0].tready),
    .probe87(axis_host_send[0].tvalid),
    .probe88(axis_host_send[1].tdata),
    .probe89(axis_host_send[1].tkeep),
    .probe90(axis_host_send[1].tlast),
    .probe91(axis_host_send[1].tready),
    .probe92(axis_host_send[1].tvalid),
    .clk(aclk)
);
`endif
