import lynxTypes::*;

/**
 * perf_fpga_axi_ctrl_parser
 * @brief Reads from/wites to the AXI Lite stream containing the benchmark data
 * 
 * @param[in] aclk Clock signal
 * @param[in] aresetn Active low reset signal
 
 * @param[in/out] axi_ctrl AXI Lite Control signal, from/to the host via PCIe and XDMA

 * @param[out] bench_ctrl Benchmark trigger to start reads/writes
 * @param[in] bench_done Number of completed reps
 * @param[in] bench_timer Benchmark timer
 * @param[out] bench_vaddr Buffer virtual address for reading/writing
 * @param[out] bench_len Buffer length (size in bytes) for reading/writing
 * @param[out] bench_pid Coyote thread ID
 * @param[out] bench_n_reps Requested number (from the user software) of read/write reps
 * @param[out] bench_n_beats Number of AXI data beats (check vfpga_top.svh and README for description)
 */
module host_networking_axi_ctrl_parser (
  input  logic                        aclk,
  input  logic                        aresetn,
  
  AXI4L.s                             axi_ctrl,

  output logic [PID_BITS-1:0]         host_networking_pid, 
  output logic [VADDR_BITS-1:0]       host_rx_buff_addr, 
  output logic [VADDR_BITS-1:0]       host_rx_buff_stride,
  output logic [VADDR_BITS-1:0]       host_rx_ring_size,
  output logic [VADDR_BITS-1:0]       host_rx_meta_addr,
  output logic [VADDR_BITS-1:0]       host_rx_meta_stride,
  input  logic [VADDR_BITS-1:0]       host_rx_ring_tail,
  output logic [VADDR_BITS-1:0]       host_rx_ring_head,
  output logic [31:0]                 host_rx_irq_coalesce
);

/////////////////////////////////////
//          CONSTANTS             //
///////////////////////////////////
localparam integer N_REGS = 2;
localparam integer ADDR_MSB = $clog2(N_REGS);
localparam integer ADDR_LSB = $clog2(AXIL_DATA_BITS/8);
localparam integer AXI_ADDR_BITS = ADDR_LSB + ADDR_MSB;

/////////////////////////////////////
//          REGISTERS             //
///////////////////////////////////
// Internal AXI registers
logic [AXI_ADDR_BITS-1:0] axi_awaddr;
logic axi_awready;
logic [AXI_ADDR_BITS-1:0] axi_araddr;
logic axi_arready;
logic [1:0] axi_bresp;
logic axi_bvalid;
logic axi_wready;
logic [AXIL_DATA_BITS-1:0] axi_rdata;
logic [1:0] axi_rresp;
logic axi_rvalid;
logic aw_en;

// Registers for holding the values read from/to be written to the AXI Lite interface
// These are synchronous but the outputs are combinatorial
logic [N_REGS-1:0][AXIL_DATA_BITS-1:0] ctrl_reg;
logic ctrl_reg_rden;
logic ctrl_reg_wren;

/////////////////////////////////////
//         REGISTER MAP           //
///////////////////////////////////

// 0 (WO)   : Buffer virtual address
localparam integer HOST_NETWORKING_PID_REG = 0;
localparam integer HOST_NETWORKING_BUFF_VADDR_REG = 1;
localparam integer HOST_NETWORKING_BUFF_STRIDE_REG = 2;
localparam integer HOST_NETWORKING_RING_SIZE_REG = 3;
localparam integer HOST_NETWORKING_META_VADDR_REG = 4;
localparam integer HOST_NETWORKING_META_STRIDE_REG = 5;
localparam integer HOST_NETWORKING_RING_TAIL_REG = 6;
localparam integer HOST_NETWORKING_RING_HEAD_REG = 7;
localparam integer HOST_NETWORKING_IRQ_COALESCE_REG = 8;

/////////////////////////////////////
//         WRITE PROCESS          //
///////////////////////////////////
// Data coming in from host to the vFPGA vie PCIe and XDMA
assign ctrl_reg_wren = axi_wready && axi_ctrl.wvalid && axi_awready && axi_ctrl.awvalid;

always_ff @(posedge aclk) begin
  if (aresetn == 1'b0) begin
    ctrl_reg <= 0;
  end
  else begin

    if(ctrl_reg_wren) begin
      case (axi_awaddr[ADDR_LSB+:ADDR_MSB])
    
        HOST_NETWORKING_PID_REG:    // Buffer virtual address
          for (int i = 0; i < (AXIL_DATA_BITS/8); i++) begin
            if(axi_ctrl.wstrb[i]) begin
              ctrl_reg[HOST_NETWORKING_PID_REG][(i*8)+:8] <= axi_ctrl.wdata[(i*8)+:8];
            end
          end

        HOST_NETWORKING_BUFF_VADDR_REG:      // Coyote Thread ID (PID)
          for (int i = 0; i < (AXIL_DATA_BITS/8); i++) begin
            if(axi_ctrl.wstrb[i]) begin
              ctrl_reg[HOST_NETWORKING_BUFF_VADDR_REG][(i*8)+:8] <= axi_ctrl.wdata[(i*8)+:8];
            end
          end

        HOST_NETWORKING_BUFF_STRIDE_REG:    // Buffer virtual address
          for (int i = 0; i < (AXIL_DATA_BITS/8); i++) begin
            if(axi_ctrl.wstrb[i]) begin
              ctrl_reg[HOST_NETWORKING_BUFF_STRIDE_REG][(i*8)+:8] <= axi_ctrl.wdata[(i*8)+:8];
            end
          end

        HOST_NETWORKING_RING_SIZE_REG:      // Coyote Thread ID (PID)
          for (int i = 0; i < (AXIL_DATA_BITS/8); i++) begin
            if(axi_ctrl.wstrb[i]) begin
              ctrl_reg[HOST_NETWORKING_RING_SIZE_REG][(i*8)+:8] <= axi_ctrl.wdata[(i*8)+:8];
            end
          end

        HOST_NETWORKING_META_VADDR_REG:    // Buffer virtual address
          for (int i = 0; i < (AXIL_DATA_BITS/8); i++) begin
            if(axi_ctrl.wstrb[i]) begin
              ctrl_reg[HOST_NETWORKING_META_VADDR_REG][(i*8)+:8] <= axi_ctrl.wdata[(i*8)+:8];
            end
          end

        HOST_NETWORKING_META_STRIDE_REG:      // Coyote Thread ID (PID)
          for (int i = 0; i < (AXIL_DATA_BITS/8); i++) begin
            if(axi_ctrl.wstrb[i]) begin
              ctrl_reg[HOST_NETWORKING_META_STRIDE_REG][(i*8)+:8] <= axi_ctrl.wdata[(i*8)+:8];
            end
          end

        HOST_NETWORKING_RING_HEAD_REG:      // Coyote Thread ID (PID)
          for (int i = 0; i < (AXIL_DATA_BITS/8); i++) begin
            if(axi_ctrl.wstrb[i]) begin
              ctrl_reg[HOST_NETWORKING_RING_HEAD_REG][(i*8)+:8] <= axi_ctrl.wdata[(i*8)+:8];
            end
          end

        HOST_NETWORKING_IRQ_COALESCE_REG:      // Coyote Thread ID (PID)
          for (int i = 0; i < (AXIL_DATA_BITS/8); i++) begin
            if(axi_ctrl.wstrb[i]) begin
              ctrl_reg[HOST_NETWORKING_IRQ_COALESCE_REG][(i*8)+:8] <= axi_ctrl.wdata[(i*8)+:8];
            end
          end

        default: ;
      endcase
    end
  end
end    

/////////////////////////////////////
//       OUTPUT ASSIGNMENT        //
///////////////////////////////////
always_comb begin
  host_rx_buff_addr             = ctrl_reg[HOST_NETWORKING_BUFF_VADDR_REG][VADDR_BITS-1:0];
  host_networking_pid           = ctrl_reg[HOST_NETWORKING_PID_REG][PID_BITS-1:0];
  host_rx_buff_stride           = ctrl_reg[HOST_NETWORKING_BUFF_STRIDE_REG][VADDR_BITS-1:0];
  host_rx_ring_size             = ctrl_reg[HOST_NETWORKING_RING_SIZE_REG][VADDR_BITS-1:0];
  host_rx_meta_addr             = ctrl_reg[HOST_NETWORKING_META_VADDR_REG][VADDR_BITS-1:0];
  host_rx_meta_stride           = ctrl_reg[HOST_NETWORKING_META_STRIDE_REG][VADDR_BITS-1:0];
  host_rx_ring_head             = ctrl_reg[HOST_NETWORKING_RING_HEAD][VADDR_BITS-1:0];
  host_rx_irq_coalesce          = ctrl_reg[HOST_NETWORKING_IRQ_COALESCE_REG][31:0];
end

/////////////////////////////////////
//       READ PROCESS              //
/////////////////////////////////////
assign ctrl_reg_rden = axi_arready & axi_ctrl.arvalid & ~axi_rvalid;

always_ff @(posedge aclk) begin
  if(aresetn == 1'b0) begin
    axi_rdata <= 0;
  end
  else begin
    if(ctrl_reg_rden) begin
      axi_rdata <= 0;

      case (axi_araddr[ADDR_LSB+:ADDR_MSB])
        HOST_NETWORKING_RING_TAIL_REG:   // Number of completions
          axi_rdata[31:0] <= host_rx_ring_tail;
        default: ;
      endcase
    end
  end 
end

/////////////////////////////////////
//     STANDARD AXI CONTROL       //
///////////////////////////////////
// NOT TO BE EDITED

// I/O
assign axi_ctrl.awready = axi_awready;
assign axi_ctrl.arready = axi_arready;
assign axi_ctrl.bresp = axi_bresp;
assign axi_ctrl.bvalid = axi_bvalid;
assign axi_ctrl.wready = axi_wready;
assign axi_ctrl.rdata = axi_rdata;
assign axi_ctrl.rresp = axi_rresp;
assign axi_ctrl.rvalid = axi_rvalid;

// awready and awaddr
always_ff @(posedge aclk) begin
  if ( aresetn == 1'b0 )
    begin
      axi_awready <= 1'b0;
      axi_awaddr <= 0;
      aw_en <= 1'b1;
    end 
  else
    begin    
      if (~axi_awready && axi_ctrl.awvalid && axi_ctrl.wvalid && aw_en)
        begin
          axi_awready <= 1'b1;
          aw_en <= 1'b0;
          axi_awaddr <= axi_ctrl.awaddr;
        end
      else if (axi_ctrl.bready && axi_bvalid)
        begin
          aw_en <= 1'b1;
          axi_awready <= 1'b0;
        end
      else           
        begin
          axi_awready <= 1'b0;
        end
    end 
end  

// arready and araddr
always_ff @(posedge aclk) begin
  if ( aresetn == 1'b0 )
    begin
      axi_arready <= 1'b0;
      axi_araddr  <= 0;
    end 
  else
    begin    
      if (~axi_arready && axi_ctrl.arvalid)
        begin
          axi_arready <= 1'b1;
          axi_araddr  <= axi_ctrl.araddr;
        end
      else
        begin
          axi_arready <= 1'b0;
        end
    end 
end    

// bvalid and bresp
always_ff @(posedge aclk) begin
  if ( aresetn == 1'b0 )
    begin
      axi_bvalid  <= 0;
      axi_bresp   <= 2'b0;
    end 
  else
    begin    
      if (axi_awready && axi_ctrl.awvalid && ~axi_bvalid && axi_wready && axi_ctrl.wvalid)
        begin
          axi_bvalid <= 1'b1;
          axi_bresp  <= 2'b0;
        end                   
      else
        begin
          if (axi_ctrl.bready && axi_bvalid) 
            begin
              axi_bvalid <= 1'b0; 
            end  
        end
    end
end

// wready
always_ff @(posedge aclk) begin
  if ( aresetn == 1'b0 )
    begin
      axi_wready <= 1'b0;
    end 
  else
    begin    
      if (~axi_wready && axi_ctrl.wvalid && axi_ctrl.awvalid && aw_en )
        begin
          axi_wready <= 1'b1;
        end
      else
        begin
          axi_wready <= 1'b0;
        end
    end 
end  

// rvalid and rresp
always_ff @(posedge aclk) begin
  if ( aresetn == 1'b0 )
    begin
      axi_rvalid <= 0;
      axi_rresp  <= 0;
    end 
  else
    begin    
      if (axi_arready && axi_ctrl.arvalid && ~axi_rvalid)
        begin
          axi_rvalid <= 1'b1;
          axi_rresp  <= 2'b0;
        end   
      else if (axi_rvalid && axi_ctrl.rready)
        begin
          axi_rvalid <= 1'b0;
        end                
    end
end    

endmodule