/**
 * This file is part of the Coyote <https://github.com/fpgasystems/Coyote>
 *
 * MIT Licence
 * Copyright (c) 2021-2025, Systems Group, ETH Zurich
 * All rights reserved.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:

 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.

 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
 */

`timescale 1ns / 1ps

import lynxTypes::*;

module tcp_notify_arb (
    // HOST 
    metaIntf.s                          s_notify,

    metaIntf.m                          m_notify_opened,
    metaIntf.m                          m_notify_recv, 

    input  logic    					aclk,    
	input  logic    					aresetn
);

metaIntf #(.STYPE(tcp_notify_t)) notify_opened (.*);
metaIntf #(.STYPE(tcp_notify_t)) notify_recv (.*);

// DP
always_comb begin
    s_notify.ready = 1'b0;

    notify_opened.valid = 1'b0;
    notify_recv.valid = 1'b0;

    if(s_notify.valid) begin
        if(s_notify.data.opened) begin
            notify_opened.valid = 1'b1;
            s_notify.ready = notify_opened.ready;
        end
        else begin
            notify_recv.valid = 1'b1;
            s_notify.ready = notify_recv.ready;
        end
    end
end

assign notify_opened.data = s_notify.data;
assign notify_recv.data = s_notify.data;

meta_reg #(.DATA_BITS($bits(tcp_notify_t))) inst_reg_0  (.aclk(aclk), .aresetn(aresetn), .s_meta(notify_opened), .m_meta(m_notify_opened));
meta_reg #(.DATA_BITS($bits(tcp_notify_t))) inst_reg_1  (.aclk(aclk), .aresetn(aresetn), .s_meta(notify_recv), .m_meta(m_notify_recv));
    
endmodule