/**
 * This file is part of the Coyote <https://github.com/fpgasystems/Coyote>
 *
 * MIT Licence
 * Copyright (c) 2021-2025, Systems Group, ETH Zurich
 * All rights reserved.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:

 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.

 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
 */

`timescale 1ns / 1ps

import lynxTypes::*;

module axis_reg_static (
	input logic 			aclk,
	input logic 			aresetn,
	
	AXI4S.s				s_axis,
	AXI4S.m 				m_axis
);

axis_register_slice_static_512 inst_reg_slice (
	.aclk(aclk),
	.aresetn(aresetn),
	.s_axis_tvalid(s_axis.tvalid),
	.s_axis_tready(s_axis.tready),
	.s_axis_tdata(s_axis.tdata),
	.s_axis_tkeep(s_axis.tkeep),
	.s_axis_tlast(s_axis.tlast),
	.m_axis_tvalid(m_axis.tvalid),
	.m_axis_tready(m_axis.tready),
	.m_axis_tdata(m_axis.tdata),
	.m_axis_tkeep(m_axis.tkeep),
	.m_axis_tlast(m_axis.tlast)
);

endmodule