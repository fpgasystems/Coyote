package simTypes;
    // --------------------------------------------------------------------------
    // CUSTOM STRUCTS
    // These are the structs to edit to adapt to any custom DUT.
    // --------------------------------------------------------------------------
    typedef struct packed {
        integer n_trs;
        integer delay;
    } c_struct_t;
    
endpackage