/**
 * This file is part of the Coyote <https://github.com/fpgasystems/Coyote>
 *
 * MIT Licence
 * Copyright (c) 2025, Systems Group, ETH Zurich
 * All rights reserved.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:

 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.

 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
 */

`timescale 1ns / 1ps

import lynxTypes::*;

/**
 * RDMA Compression Engine
 *
 * This module implements a framework for data compression on RDMA traffic.
 * The compression operates on 512-bit AXI streams at 250 MHz to support 100G line rate.
 *
 * Design Features:
 * - Zero backpressure: always accepts data when ready
 * - Pipelined design for high throughput
 * - Metadata preservation: tid, tlast, tkeep signals are maintained
 * - Extensible framework for implementing compression algorithms
 *
 * Current Implementation:
 * - Passthrough mode with compression statistics tracking
 * - Detects zero patterns for compression ratio estimation
 * - Ready for extension with actual compression algorithms (RLE, LZ77, Snappy, etc.)
 *
 * To implement actual compression:
 * - Replace the passthrough logic in Stage 1 with compression algorithm
 * - Modify output format to include compressed data and metadata
 * - Ensure decompression module implements the reverse transformation
 */
module rdma_compression_engine (
    input  logic        aclk,
    input  logic        aresetn,
    
    // Input AXI Stream (from host/network)
    AXI4SR.s            axis_in,
    
    // Output AXI Stream (to network/host, compressed)
    AXI4SR.m            axis_out
);

    // Pipeline stages for maintaining throughput
    localparam int PIPELINE_DEPTH = 2;
    
    // Internal pipeline signals
    AXI4SR axis_pipe[PIPELINE_DEPTH+1]();
    
    // Stage 0: Input buffer/register
    axisr_reg inst_input_reg (
        .aclk(aclk),
        .aresetn(aresetn),
        .s_axis(axis_in),
        .m_axis(axis_pipe[0])
    );
    
    // Stage 1: Compression logic
    // For this demonstration, we implement a passthrough with compression statistics
    // In a real implementation, this would contain the actual compression algorithm
    logic [AXI_DATA_BITS-1:0] compressed_data;
    logic compressed_valid;
    logic [63:0] compression_ratio_counter;
    
    always_ff @(posedge aclk) begin
        if (~aresetn) begin
            compressed_valid <= 1'b0;
            compression_ratio_counter <= 64'h0;
        end else begin
            compressed_valid <= axis_pipe[0].tvalid;
            compressed_data <= axis_pipe[0].tdata;
            
            // Simple compression: detect zero patterns
            // In production, this would be a more sophisticated algorithm
            if (axis_pipe[0].tvalid && axis_pipe[0].tready) begin
                // Check if data is all zeros (highly compressible)
                if (axis_pipe[0].tdata == '0) begin
                    compression_ratio_counter <= compression_ratio_counter + 1;
                end
            end
        end
    end
    
    // Assign compressed data to pipeline stage 1
    assign axis_pipe[1].tdata = compressed_data;
    assign axis_pipe[1].tvalid = compressed_valid;
    assign axis_pipe[1].tkeep = axis_pipe[0].tkeep;
    assign axis_pipe[1].tlast = axis_pipe[0].tlast;
    assign axis_pipe[1].tid = axis_pipe[0].tid;
    assign axis_pipe[0].tready = axis_pipe[1].tready;
    
    // Stage 2: Output buffer/register
    axisr_reg inst_output_reg (
        .aclk(aclk),
        .aresetn(aresetn),
        .s_axis(axis_pipe[1]),
        .m_axis(axis_out)
    );

endmodule

/**
 * RDMA Decompression Engine
 *
 * This module implements a framework for data decompression on RDMA traffic.
 * It operates on 512-bit AXI streams at 250 MHz to support 100G line rate.
 *
 * Design Features:
 * - Zero backpressure: always accepts data when ready
 * - Pipelined design for high throughput
 * - Metadata preservation: tid, tlast, tkeep signals are maintained
 * - Extensible framework for implementing decompression algorithms
 *
 * Current Implementation:
 * - Passthrough mode with decompression statistics tracking
 * - Symmetric to the compression engine's passthrough mode
 * - Ready for extension with actual decompression algorithms
 *
 * To implement actual decompression:
 * - Replace the passthrough logic in Stage 1 with decompression algorithm
 * - Must match the compression format implemented in rdma_compression_engine
 * - Parse compressed data and metadata to reconstruct original data
 */
module rdma_decompression_engine (
    input  logic        aclk,
    input  logic        aresetn,
    
    // Input AXI Stream (compressed data from network/host)
    AXI4SR.s            axis_in,
    
    // Output AXI Stream (decompressed data to host/network)
    AXI4SR.m            axis_out
);

    // Pipeline stages for maintaining throughput
    localparam int PIPELINE_DEPTH = 2;
    
    // Internal pipeline signals
    AXI4SR axis_pipe[PIPELINE_DEPTH+1]();
    
    // Stage 0: Input buffer/register
    axisr_reg inst_input_reg_decomp (
        .aclk(aclk),
        .aresetn(aresetn),
        .s_axis(axis_in),
        .m_axis(axis_pipe[0])
    );
    
    // Stage 1: Decompression logic
    logic [AXI_DATA_BITS-1:0] decompressed_data;
    logic decompressed_valid;
    logic [63:0] decompression_counter;
    
    always_ff @(posedge aclk) begin
        if (~aresetn) begin
            decompressed_valid <= 1'b0;
            decompression_counter <= 64'h0;
        end else begin
            decompressed_valid <= axis_pipe[0].tvalid;
            decompressed_data <= axis_pipe[0].tdata;
            
            // Decompression logic
            // In production, this would reverse the compression algorithm
            if (axis_pipe[0].tvalid && axis_pipe[0].tready) begin
                decompression_counter <= decompression_counter + 1;
            end
        end
    end
    
    // Assign decompressed data to pipeline stage 1
    assign axis_pipe[1].tdata = decompressed_data;
    assign axis_pipe[1].tvalid = decompressed_valid;
    assign axis_pipe[1].tkeep = axis_pipe[0].tkeep;
    assign axis_pipe[1].tlast = axis_pipe[0].tlast;
    assign axis_pipe[1].tid = axis_pipe[0].tid;
    assign axis_pipe[0].tready = axis_pipe[1].tready;
    
    // Stage 2: Output buffer/register
    axisr_reg inst_output_reg_decomp (
        .aclk(aclk),
        .aresetn(aresetn),
        .s_axis(axis_pipe[1]),
        .m_axis(axis_out)
    );

endmodule
