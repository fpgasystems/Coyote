/**
 * This file is part of the Coyote <https://github.com/fpgasystems/Coyote>
 *
 * MIT Licence
 * Copyright (c) 2021-2025, Systems Group, ETH Zurich
 * All rights reserved.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:

 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.

 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
 */

`timescale 1ns / 1ps

import lynxTypes::*;

module dcpl_select #(
    parameter integer                       N_STAGES = 1,
    parameter integer                       N_DCPL = N_REGIONS
) (
    input  logic                            aclk,
    input  logic                            aresetn,
    
    input  logic [N_DCPL-1:0]               decouple_sw,
    output logic [N_DCPL-1:0]               decouple
);  

    logic [N_STAGES:0][N_DCPL-1:0] decouple_out;

    // I/O
    assign decouple_out[0] = decouple_sw;
    assign decouple = decouple_out[N_STAGES];

    // Reg
    always_ff @(posedge aclk) begin
        if(~aresetn) begin
            for(int i = 1; i <= N_STAGES; i++) begin
                decouple_out[i] <= 0;
            end
        end
        else begin
            for(int i = 1; i <= N_STAGES; i++) begin
                decouple_out[i] <= decouple_out[i-1];
            end
        end
    end
    
endmodule
