/*
    Copyright (c) 2022 ETH Zurich.
    All rights reserved.

    This file is distributed under the terms in the attached LICENSE file.
    If you do not find this file, copies can be found by writing to:
    ETH Zurich D-INFK, Stampfenbachstrasse 114, CH-8092 Zurich. Attn: Systems Group
*/

/*

	The link_state_machine module maintains the link state. It operates in three different phases:
	1- Init Phase: in this phase the link state machine exchanges init requests and acknowledgement with its
	   partner on the other side of the link.
	2- Run phase: int this phase the link state machine allow the exchange od data/credit blocks.
	3- Error handling phase: in this phase the link state machine react for errors detected while receiving blocks
	   or errors detected by its partner.


	When first reset, the state machine is in the IREQ state, the state machine responds
	to a valid sync block and error messages. If none, it stays in its current state.

	States:

	Init Phase: this phase covers the IREQ and IACK states. The link state machine enters this phase on
	            a global reset (rst_n signal active low), when the partner on the link request link reinitialization,
	            or when the link state machine receives csr init request.  The Init Phase starts with the IREQ
	            state, and on receiving init ack from the partner, it moves to the IACK state, until the partner
	            stop acknowledging and generating init requests, then the link state machine moves to the RUN state.

	Run Phase: This phase covers the RUN state. In this phase, the link state machine monitors errors and partner
			   init or retry requests. If no such signal detected, data blocks are generated or IDLE blocks if there
			   is no data.

	Error phase: This phase covers three states: RREQ, RACK, REPLAY. In this phase there are two behaviors
				for the link state machine, first if it detects an error in the received blocks then it enters the
				RREQ state to generate a retry request, once the partner acknowledge it, it moves to the RACK state
				until the partner stops acknowledging requests then it moves back to the RUN state.
				The second behavior is triggered by retry requests generated by the partner, then it moves to the
				RACK state to acknowledge the retry requests, once the partner receives the acknowledgement it moves
				to the REPLAY state to resend latest blocks stored in the REPLAY buffer. Once it is done, it moves
				back to the RUN state. The comlexity of this phase comes from the fact that these two behaviors
				can overlap in any of the thre states.

	IREQ:
		Generate SYNC blocks with Req[1:0] = 01
		if receives InitAck then it moves to IACK state
		output: {7x64b0}{ 3'b110, 1'b0, 6'b0, 2'b01, 12'b0, 8'b0, 8'b0, CRC}

	IACK:
		On entrance to this state it starts generating Synch blocks with Req[1:0] = 00
		When it receives an InitReq then it asserts InitAck
		When both received InitAck or InitReq are deasserted, it moves to the RUN state
		Output: on entrance: {7x64b0} { 3'b110, 1'b0, 6'b0, 2'b00, 12'b0, 7'b0, 7'b0, CRC}
				on InitReq:  {7x64b0} { 3'b110, 1'b1, 6'b0, 2'b00, 12'b0, 7'b0, 7'b0, CRC}
	RUN:
		In this state Generate block unit is allowed to receive data and send IDLE blocks
		if no data or credit available.

		Immediatelly on entering this state, credit blocks are generated without data
		to return credit to the partner.

		If an error is detected in the received blocks, the generate block stops transmiting data
		and enters the RREQ state.

		If a RetryReq received in the RX then it issues a RetryAck and enters RACK state

	RREQ:
		In this states it generates SYNC blocks with Req[1:0] = 11, until it receives RetryAck
		then it deasserts the RetryReq and goes to RACK state.



*/


import block_types::*;


module link_state_machine (
	input   wire 						clk,                        // Clock
	input   wire 						rst_n,                      // Asynchronous reset active low

	//------------  Inputs from the Block RX Path ------------//
	input   SyncBlock_t   				rx_sync_block,              // Sync Block from RLK
	input   wire 						rx_sync_block_valid,
	input   wire                        rx_blk_received,         	// A valid data block received
	input   wire 						rx_blk_error,               // CRC error detected

	//--------------- Input Data from Arbiter ----------------//
	input   DataBlock_t                 arb_data_block,
	input   wire 						arb_data_block_valid,
	output  wire 						arb_data_block_ready,

	//----------------- Credits to Return --------------------//
	input   wire [12:0]                 rx_vc_fifo_pop,       // if a bit is 1 => 8 words poped from the VC RX FIFO

	input   wire 						csr_init,
	output  wire 						link_up,
	output  wire [5:0]     				out_link_state,

	// Output Block
	output  wire [BLOCK_WIDTH-1:0] 		tx_block_out,
	input   wire 						tx_block_out_ready,

	//------------------- Debug Output ----------------------//
	output  wire  [63:0] 				debug_counters,
	output  wire  [95:0] 				debug_counters2,
	output  reg   [5:0] 				blk_trx_state

);

Block_t 				tx_block_out_t;

// {B5: Replay bit, B4:B3: Retry bit, B2: Run bit, B1: Init bit, B0 Request bit}

localparam   [5:0]    IREQ   = 6'b000001,
					  IACK   = 6'b000010,
					  RUN    = 6'b000100,
					  RREQ   = 6'b001000,
					  RACK   = 6'b010000,
					  REPLAY = 6'b100000;


reg                                 rx_sync_block_valid_d1;
SyncBlock_t                      	rx_sync_block_d1;
SyncBlock_t                      	tx_sync_block_w1;

DataBlock_t							data_block;
DataBlock_t							replay_block;
DataBlock_t							idle_block;
DataBlock_t						 	credit_block;

DataBlock_t                         replay_mem_din;
wire 								replay_mem_we;
reg     [7:0] 						replay_mem_waddr;
wire 								replay_mem_re;
reg     [7:0] 						replay_mem_raddr;
reg     [7:0] 						next_replay_mem_raddr;


SyncBlock_t 					 	sync_block;

reg 							 	rx_init_req;
reg 								rx_retry_req;
reg 							 	rx_init_ack;
reg 							 	rx_retry_ack;
reg 	[7:0]					  	retry_seq;

reg 	[7:0]					 	tx_seq;
wire  	[7:0]					 	tx_seq_minus_1;
reg     [5:0]					  	link_state;
reg     [5:0]					  	link_state_sending;
reg     [5:0]					  	next_link_state;
reg     [5:0]					  	prev_link_state;

reg 								rack_error;
reg 							 	tlk_blk_retry;
reg 								replay_needed;
reg 	[23:0] 						rreq_timer;

reg 								next_tlk_blk_retry;
reg 	[23:0]						next_rreq_timer;

// NOT IMPLEMENTED YET
wire    [7:0] 						retry_ptr;
wire 								return_ack;
reg     [6:0] 						ack_cnt;
reg 								last_replay;
wire 								last_replay_w;
wire 								last_replay_sent;
DataBlock_t			 				replay_mem_block;
reg     [7:0] 						rx_seq;

//
reg   	[3:0] 						ireq_iack_moves;
reg   	[3:0] 						iack_run_moves;
reg   	[3:0] 						iack_rreq_moves;
reg   	[3:0] 						run_rreq_moves;
reg   	[3:0] 						run_rack_moves;
reg   	[3:0] 						run_ireq_moves;

reg   	[3:0] 						rreq_rack_moves;
reg   	[3:0] 						rreq_ireq_moves;
reg   	[3:0] 						rack_ireq_moves;
reg   	[3:0] 						rack_run_moves;
reg   	[3:0] 						rack_rreq_moves;
reg   	[3:0] 						rack_replay_moves;

reg   	[3:0] 						replay_ireq_moves;
reg   	[3:0] 						replay_rreq_moves;
reg   	[3:0] 						replay_run_moves;
reg   	[3:0] 						replay_rack_moves;

reg   	[15:0] 						rx_retry_req_rises;
reg   	[15:0] 						rx_retry_req_falls;
reg   	[15:0] 						rx_retry_ack_rises;
reg   	[15:0] 						rx_retry_ack_falls;

reg  	[8:0]    					vc_credit[12:0];
wire 	[12:0]   					vc_credit_to_return;
reg  	[12:0]   					vc_credit_dec;
reg  		  						high_first;
reg  	[7:0]    					credits_to_return;
reg 								block_type;
wire 		  						credit_tx_ready;

reg     [15:0]                      replay_blocks_count;
reg     [11:0]                      cred_blocks_count;
reg     [3:0]                       retry_req_sent;

//////////////////////////////////////////////////////////////////////////
//////////////////////         Debug Counters         ////////////////////
//////////////////////////////////////////////////////////////////////////

assign  debug_counters = {replay_rack_moves, replay_run_moves, replay_rreq_moves, replay_ireq_moves,
						  rack_replay_moves, rack_rreq_moves, rack_run_moves, rack_ireq_moves,
						  rreq_ireq_moves, rreq_rack_moves, run_ireq_moves, run_rack_moves,
						  run_rreq_moves, iack_rreq_moves, iack_run_moves, ireq_iack_moves};

assign debug_counters2 = {retry_req_sent, cred_blocks_count, replay_blocks_count, rx_retry_req_rises, rx_retry_req_falls, rx_retry_ack_rises, rx_retry_ack_falls};

always@(posedge clk) begin
	if(~rst_n) begin
		ireq_iack_moves  <= 4'h0;
		iack_run_moves   <= 4'h0;
		iack_rreq_moves  <= 4'h0;
		run_ireq_moves   <= 4'h0;
		run_rreq_moves   <= 4'h0;
		run_rack_moves   <= 4'h0;
		rreq_rack_moves  <= 4'h0;
		rreq_ireq_moves  <= 4'h0;
		rack_run_moves   <= 4'h0;
		rack_ireq_moves  <= 4'h0;
		rack_replay_moves<= 4'h0;
		rack_rreq_moves  <= 4'h0;
		replay_ireq_moves<= 4'h0;
		replay_rreq_moves<= 4'h0;
		replay_run_moves <= 4'h0;
		replay_rack_moves<= 4'h0;

		blk_trx_state    <= 6'b0;

		prev_link_state  <= 6'b0;

		rx_retry_req_rises <= 16'b0;
		rx_retry_req_falls <= 16'b0;

		rx_retry_ack_rises <= 16'b0;
		rx_retry_ack_falls <= 16'b0;

	end
	else begin
		prev_link_state  <= link_state;
		blk_trx_state    <= link_state;


		ireq_iack_moves <= 	(ireq_iack_moves == 4'hF)? ireq_iack_moves :
							(prev_link_state[0] & link_state[1])? ireq_iack_moves + 1'b1 : ireq_iack_moves;

		iack_run_moves  <= 	(iack_run_moves == 4'hF)? iack_run_moves :
							(prev_link_state[1] & link_state[2])? iack_run_moves + 1'b1  : iack_run_moves;

		iack_rreq_moves <= 	(iack_rreq_moves == 4'hF)? iack_rreq_moves :
							(prev_link_state[1] & link_state[3])? iack_rreq_moves + 1'b1 : iack_rreq_moves;

		run_ireq_moves  <= 	(run_ireq_moves == 4'hF)? run_ireq_moves :
							(prev_link_state[2] & link_state[0])? run_ireq_moves + 1'b1 : run_ireq_moves;

		run_rreq_moves  <= 	(run_rreq_moves == 4'hF)? run_rreq_moves :
							(prev_link_state[2] & link_state[3])? run_rreq_moves + 1'b1 : run_rreq_moves;

		run_rack_moves  <= 	(run_rack_moves == 4'hF)? run_rack_moves :
							(prev_link_state[2] & link_state[4])? run_rack_moves + 1'b1 : run_rack_moves;

		rreq_rack_moves <= 	(rreq_rack_moves == 4'hF)? rreq_rack_moves :
							(prev_link_state[3] & link_state[4])? rreq_rack_moves + 1'b1 : rreq_rack_moves;

		rreq_ireq_moves <= 	(rreq_ireq_moves == 4'hF)? rreq_ireq_moves :
							(prev_link_state[3] & link_state[0])? rreq_ireq_moves + 1'b1 : rreq_ireq_moves;

		rack_run_moves  <= 	(rack_run_moves == 4'hF)? rack_run_moves :
							(prev_link_state[4] & link_state[2])? rack_run_moves + 1'b1 : rack_run_moves;

		rack_ireq_moves <= 	(rack_ireq_moves == 4'hF)? rack_ireq_moves :
							(prev_link_state[4] & link_state[0])? rack_ireq_moves + 1'b1 : rack_ireq_moves;

		rack_replay_moves<= (rack_replay_moves == 4'hF)? rack_replay_moves :
							(prev_link_state[4] & link_state[5])? rack_replay_moves + 1'b1 : rack_replay_moves;

		rack_rreq_moves <= 	(rack_rreq_moves == 4'hF)? rack_rreq_moves :
							(prev_link_state[4] & link_state[3])? rack_rreq_moves + 1'b1 : rack_rreq_moves;

		replay_ireq_moves<= (replay_ireq_moves == 4'hF)? replay_ireq_moves :
							(prev_link_state[5] & link_state[0])? replay_ireq_moves + 1'b1 : replay_ireq_moves;

		replay_rreq_moves<= (replay_rreq_moves == 4'hF)? replay_rreq_moves :
							(prev_link_state[5] & link_state[3])? replay_rreq_moves + 1'b1 : replay_rreq_moves;

		replay_run_moves <= (replay_run_moves == 4'hF)? replay_run_moves :
							(prev_link_state[5] & link_state[2])? replay_run_moves + 1'b1 : replay_run_moves;

		replay_rack_moves<= (replay_rack_moves == 4'hF)? replay_rack_moves :
							(prev_link_state[5] & link_state[4])? replay_rack_moves + 1'b1 : replay_rack_moves;


		//
		if(rx_sync_block_valid) begin

			rx_retry_req_rises <= (rx_sync_block.Req[1]  && rx_sync_block.Req[0] && !rx_retry_req)? rx_retry_req_rises + 1'b1 : rx_retry_req_rises;
			rx_retry_req_falls <= (!(rx_sync_block.Req[1]  && rx_sync_block.Req[0]) && rx_retry_req)? rx_retry_req_falls + 1'b1 : rx_retry_req_falls;

			rx_retry_ack_rises <= (rx_sync_block.Req[1]  && rx_sync_block.Ack && !rx_retry_ack)? rx_retry_req_rises + 1'b1 : rx_retry_req_rises;
			rx_retry_ack_falls <= (!(rx_sync_block.Req[1]  && rx_sync_block.Ack) && rx_retry_ack)? rx_retry_req_falls + 1'b1 : rx_retry_req_falls;
		end

	end
end

//////////////////////////////////////////////////////////////////////////
//////////////////////       Decode Sync Block        ////////////////////
//////////////////////////////////////////////////////////////////////////

// Decode Received Sync Block logic

always@(posedge clk) begin
	if(~rst_n) begin
		rx_sync_block_d1       	<= 0;
		rx_sync_block_valid_d1 	<= 1'b0;

		rx_init_ack 		 	<= 0;
		rx_init_req  			<= 0;
		rx_retry_req 			<= 0;
		rx_retry_ack 			<= 0;

		retry_seq    			<= 0;
	end
	else begin
		rx_sync_block_d1       <= rx_sync_block;
		rx_sync_block_valid_d1 <= rx_sync_block_valid;



		if(rx_sync_block_valid) begin
			rx_init_ack  <= (!rx_sync_block.Req[1] && rx_sync_block.Ack);
			rx_init_req  <= (!rx_sync_block.Req[1] && rx_sync_block.Req[0]);
			rx_retry_req <= (rx_sync_block.Req[1]  && rx_sync_block.Req[0]);
			rx_retry_ack <= (rx_sync_block.Req[1]  && rx_sync_block.Ack);

			retry_seq    <= rx_sync_block.RxSEQ;
		end
	end
end

//////////////////////////////////////////////////////////////////////////
//////////////////////      Block Acknowledgement     ////////////////////
//////////////////////////////////////////////////////////////////////////

assign return_ack = |ack_cnt[6:3];

always@(posedge clk) begin
	if(~rst_n) begin
		ack_cnt <= 7'b0;
	end
	else begin
		if(link_state[0] | link_state[1] | link_state[3] | link_state[4]) begin
			ack_cnt <= 7'b0;
		end
		else if(link_state[2] | link_state[5]) begin   // run or replay state
			if(rx_blk_received) begin
				if(tx_block_out_ready && return_ack) begin
					ack_cnt <= ack_cnt - 7'd7;
				end
				else begin
					ack_cnt <= ack_cnt + 7'd1;
				end
			end
			else if(tx_block_out_ready && return_ack) begin
				ack_cnt <= ack_cnt - 7'd8;
			end
		end
	end
end

//////////////////////////////////////////////////////////////////////////
//////////////////////          Link State            ////////////////////
//////////////////////////////////////////////////////////////////////////

assign link_up = link_state == RUN || link_state == RACK || link_state == RREQ || link_state == REPLAY;
assign out_link_state = link_state;

always@(posedge clk) begin
	if(~rst_n) begin
		link_state    <= IREQ;
        rreq_timer    <= 0;
        tlk_blk_retry <= 1'b0;

        rack_error    <= 1'b0;

        replay_needed <= 1'b0;
	end
	else begin
		link_state    <= next_link_state;
		rreq_timer    <= next_rreq_timer;
		tlk_blk_retry <= next_tlk_blk_retry;

		replay_needed <= tx_seq != retry_seq;

		if(link_state[2]) begin
			rack_error <= 1'b0;
		end
		else if(link_state[4] && rx_blk_error && !rx_init_req && !rx_retry_req) begin
			rack_error <= rx_blk_error || rack_error;
		end
	end
end

always@(*) begin
	next_link_state           = link_state;
	next_tlk_blk_retry        = 1'b0;

	//
	next_rreq_timer           = rreq_timer;

	// Output Sync Block fields
	sync_block.Type   = BTYPE_SYNC;
	sync_block.Zeros  = 6'b0;
	sync_block.Zeros2 = 12'b0;
	sync_block.Crc24  = 24'b0;
	sync_block.TxSEQ  = 8'b0;
	sync_block.RxSEQ  = 8'b0;
	sync_block.Req    = 2'b00;
	sync_block.Ack    = 1'b0;

	case (link_state)
		/* If it receives InitAck then it moves to IACK state */
		IREQ: begin
			if(rx_init_ack) begin
				next_link_state = IACK;
			end

			// Sync block fields to set in this state: send init requst, acknowledge received init requests
			sync_block.Req = 2'b01;
			sync_block.Ack = rx_init_req;

			//
			next_rreq_timer = 0;
		end
		/* If it receives an error on the RX then it moves to RREQ,
		   If both init_ack and init_req are deasserted in the RLK then we
		   move to the RUN state.
		*/
		IACK: begin
            if(rx_init_ack || rx_init_req || csr_init) begin
				next_link_state = IACK;
			end
            else if(rx_blk_error) begin
				next_link_state = RREQ;
			end
			else if(~rx_init_ack && ~rx_init_req && rx_sync_block_valid_d1) begin
				next_link_state = RUN;
			end

			// Sync block fields to set in this state: only acknowledge received init requests
			sync_block.Ack = rx_init_req;

			//
			next_rreq_timer = 0;
		end
		/* If it receives init_req from the RLK it goes back to the initial state
		   if an error is detected in the RLK received blocks then we switch to
		   the Retry Requests State (RREQ). If a Retry Request is received in the RLK
		   then we move to RACK state
		*/
		RUN: begin
			if(rx_init_req || csr_init) begin
				next_link_state = IREQ;
			end
			else if(rx_blk_error || rack_error) begin
				next_link_state = RREQ;
			end
			else if(rx_retry_req) begin
				next_link_state = RACK;
			end

			//
			next_tlk_blk_retry = rx_retry_req && replay_needed;

			//
			next_rreq_timer = 0;
		end
		/*  If it receives init_req from the RLK it goes back to the initial state
		   if an error is detected in the RLK received blocks then we stay in this state.
		   If it receives retry_ack from RLK then it moves to RACK state.
		*/
		RREQ: begin
			if(rx_init_req || csr_init) begin
				next_link_state = IREQ;
			end
			else if(rx_blk_error) begin
				next_link_state = RREQ;
			end
			else if(rx_retry_ack) begin
				next_link_state = RACK;
			end

			//
			next_tlk_blk_retry = replay_needed;

			//
			if(rx_blk_error) begin
				next_rreq_timer = 0;
			end
			else if(tx_block_out_ready) begin
                if (rreq_timer != 24'hFFFFFF) begin
				    next_rreq_timer = rreq_timer + 1'b1;
				end else begin
    				next_link_state = IREQ;
				end
			end

			// generate retry request, acknowledge retry requests set retry ptr
			sync_block.Req   = 2'b11;
			sync_block.Ack   = rx_retry_req;
			sync_block.TxSEQ = retry_ptr;
			sync_block.RxSEQ = rx_seq;
		end
		/*  If it receives init_req from the RLK it goes back to the initial state
		*/
		RACK: begin
			if(rx_init_req || csr_init) begin
				next_link_state = IREQ;
			end
			else if((rx_retry_req || rx_retry_ack)) begin
				next_link_state = RACK;
			end
			else if(rx_blk_error) begin
				next_link_state = RREQ;
			end
			else if(tlk_blk_retry) begin
				next_link_state = REPLAY;
			end
            else if (!rx_retry_ack && rx_sync_block_valid_d1) begin
                 next_link_state = RUN;
            end

            //
            next_tlk_blk_retry = replay_needed;

			//
			next_rreq_timer = 0;

            // generate retry request, acknowledge retry requests
			sync_block.Req   = 2'b10;
			sync_block.Ack   = rx_retry_req;
			sync_block.TxSEQ = retry_ptr;
			sync_block.RxSEQ = rx_seq;
		end

		REPLAY: begin
			if(rx_init_req || csr_init) begin
				next_link_state = IREQ;
			end
            else if (rx_blk_error) begin
                next_link_state = RREQ;
            end
            else if(rx_retry_req) begin
            	next_link_state = RACK;
            end
            else if (last_replay_sent) begin
                next_link_state = RUN;
            end
            //
            next_tlk_blk_retry = !last_replay_sent;
		end
		default: begin
			next_link_state    = IREQ;
			next_tlk_blk_retry = 1'b0;
		end
	endcase
end


//////////////////////////////////////////////////////////////////////////
//////////////////////    Compose Valid Data Block     ///////////////////
//////////////////////////////////////////////////////////////////////////
// append acknowledgement and credits to data block

assign arb_data_block_ready = link_state[2] && tx_block_out_ready;

assign data_block = '{Data:    arb_data_block.Data,
					  Type:    ((block_type)? BTYPE_HI : BTYPE_LO),
                      Ack:     return_ack,
                      Credits: credits_to_return,
                      Vcs:     arb_data_block.Vcs,
                      Crc24:   24'b0 };

//////////////////////////////////////////////////////////////////////////
////////////////////////    Compose Credit Block     /////////////////////
//////////////////////////////////////////////////////////////////////////
// append acknowledgement and credits

assign credit_block = '{Data:    {64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0},
					    Type:    ((block_type)? BTYPE_HI : BTYPE_LO),
                        Ack:     return_ack,
                        Credits: credits_to_return,
                        Vcs:     {4'hF, 4'hF, 4'hF, 4'hF, 4'hF, 4'hF, 4'hF},
                        Crc24:   24'b0 };

assign credit_tx_ready = link_state[2] && tx_block_out_ready;
//////////////////////////////////////////////////////////////////////////
//////////////////////    Compose Replay Data Block     //////////////////
//////////////////////////////////////////////////////////////////////////
// append acknowledgement replay block

assign replay_block = '{Data:    replay_mem_block.Data,
					    Type:    replay_mem_block.Type,
                        Ack:     return_ack,
                        Credits: replay_mem_block.Credits,
                        Vcs:     replay_mem_block.Vcs,
                        Crc24:   24'b0 };

//////////////////////////////////////////////////////////////////////////
/////////////////////////    Compose Idle Block     //////////////////////
//////////////////////////////////////////////////////////////////////////
// append acknowledgement

assign idle_block   = '{Data:    {64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0},
					    Type:    BTYPE_IDLE,
                        Ack:     return_ack,
                        Credits: 8'b0,
                        Vcs:     {4'hF, 4'hF, 4'hF, 4'hF, 4'hF, 4'hF, 4'hF},
                        Crc24:   24'b0 };

//////////////////////////////////////////////////////////////////////////
/////////////////////////    Select Output Block     /////////////////////
//////////////////////////////////////////////////////////////////////////

always@(posedge clk) begin
	if(~rst_n) begin
		tx_block_out_t <= '{Data:          {64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0},
					  	  custom_fields: {idle_block.Type, idle_block.Ack, 8'h00, tx_seq, rx_seq, 12'h000},
					      Crc24:         24'b0};

		tx_seq             <= 8'b0;
		link_state_sending <= IREQ;
	end
	else if(tx_block_out_ready) begin
		link_state_sending <= link_state;
		case (link_state)
			RUN: begin
				if(arb_data_block_valid) begin
					tx_block_out_t <= '{Data:         data_block.Data,
					  	  			  custom_fields: {data_block.Type, data_block.Ack, data_block.Credits, data_block.Vcs},
					      			  Crc24:         24'b0};

					tx_seq       <= tx_seq + 1'b1;
				end
				else if(|credits_to_return) begin
					tx_block_out_t <= '{Data:         {64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0},
					  	  			  custom_fields: {credit_block.Type, credit_block.Ack, credit_block.Credits, 28'hFFFFFFF},
					      			  Crc24:         24'b0};

					tx_seq       <= tx_seq + 1'b1;
				end
				else begin
					tx_block_out_t <= '{Data:         {64'b0, 4'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0},
					  	  			  custom_fields: {idle_block.Type, idle_block.Ack, 8'h00, retry_ptr, rx_seq, 12'h000},
					      			  Crc24:         24'b0};
				end
			end
			REPLAY: begin
				tx_block_out_t <= '{Data:         replay_block.Data,
					  	  	      custom_fields: {replay_block.Type, replay_block.Ack, replay_block.Credits, replay_block.Vcs},
					      		  Crc24:         24'b0};
			end
			IREQ, IACK, RREQ, RACK: begin
				tx_block_out_t <= '{Data:         {64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0},
					  	  	      custom_fields: {sync_block.Type, sync_block.Ack, sync_block.Zeros, sync_block.Req, sync_block.TxSEQ, sync_block.RxSEQ, sync_block.Zeros2},
					      		  Crc24:         24'b0};

				tx_seq       <= (link_state[0] | link_state[1])? 8'b0 : tx_seq;
			end
			default : begin
				tx_block_out_t <= '{Data:          {64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0, 64'b0},
					  	  		  custom_fields: {idle_block.Type, idle_block.Ack, 8'h00, retry_ptr, rx_seq, 12'h000},
					      		  Crc24:         24'b0};
				tx_seq       <= 8'b0;
			end
		endcase
	end
end

assign tx_block_out = {tx_block_out_t.Data,
                      tx_block_out_t.custom_fields,
                      tx_block_out_t.Crc24};

assign tx_seq_minus_1   = tx_seq - 1'b1;
////////////////////////////////////////////////////

always@(posedge clk) begin
	if(~rst_n) begin
		rx_seq              <= 0;
	//	retry_ptr           <= 0;
	end
	else begin
		// rx_seq
		if( |link_state[1:0]) begin
			rx_seq <= 0;
		end
		else if(rx_blk_received) begin
			rx_seq <= rx_seq + 1'b1;
		end
		/*// retry_ptr
		if(link_state[0] | link_state[1]) begin
			retry_ptr <= 0;
		end
		else if(link_state[4]) begin
			retry_ptr <= retry_seq;
		end
		else if(link_state[5] && !last_replay && tx_block_out_ready) begin
			retry_ptr <= retry_ptr + 1'b1;
		end*/
	end
end

////////////////////////////////////////////////////
// DEBUG COUNTERS
always@(posedge clk) begin
	if(~rst_n) begin
		replay_blocks_count <= 0;
		cred_blocks_count   <= 0;
		retry_req_sent      <= 0;
	end
	else begin
		//
		if(tx_block_out_ready && link_state[5] && (replay_blocks_count != 16'hFFFF)) begin
			replay_blocks_count <= replay_blocks_count + 1'b1;
		end
		//
		if(credit_tx_ready && (|credits_to_return) && (cred_blocks_count != 12'hFFF)) begin
			cred_blocks_count <= cred_blocks_count + 1'b1;
		end
		//
		if(tx_block_out_ready &&  (&(tx_block_out_t.custom_fields[29:28])) && (retry_req_sent != 4'hF) &&  (tx_block_out_t.custom_fields[38:37] != 2'b10) ) begin
			retry_req_sent <= retry_req_sent + 1'b1;
		end
		//

	end
end

//////////////////////////////////////////////////////////////////////////
/////////////////////////    VC Returned Credit      /////////////////////
//////////////////////////////////////////////////////////////////////////

// vc_credit_dec: decrement credit counters whenever a credit return word is sent.
always@(*) begin
	vc_credit_dec = 13'b0;

	if(credit_tx_ready) begin
		if(high_first) begin
			if(|vc_credit_to_return[12:8]) begin
				vc_credit_dec = {vc_credit_to_return[12:8], 8'h00};
			end
			else begin
				vc_credit_dec = {5'b00000, vc_credit_to_return[7:0]};
			end
		end
		else begin
			if(|vc_credit_to_return[7:0]) begin
				vc_credit_dec = {5'b00000, vc_credit_to_return[7:0]};
			end
			else begin
				vc_credit_dec = {vc_credit_to_return[12:8], 8'h00};
			end
		end
	end
end

// high_first: flag bit to arbitrate between high and low channels.
// credits_to_return: credits word to be returned.
always@(posedge clk) begin
	if(~rst_n) begin
		high_first  	  <= 1'b0;
		credits_to_return <= 8'b0;
		block_type        <= 1'b0;
	end
	else if(credit_tx_ready) begin
		if(high_first) begin
			if(|vc_credit_to_return[12:8]) begin
				high_first        <= 1'b0;
				credits_to_return <= {3'b000, vc_credit_to_return[12:8]};
				block_type        <= 1'b1;
			end
			else begin
				credits_to_return <= vc_credit_to_return[7:0];
				block_type        <= 1'b0;
			end
		end
		else begin
			if(|vc_credit_to_return[7:0]) begin
				high_first        <= 1'b1;
				credits_to_return <= vc_credit_to_return[7:0];
				block_type        <= 1'b0;
			end
			else begin
				credits_to_return <= {3'b000, vc_credit_to_return[12:8]};
				block_type        <= 1'b1;
			end
		end
	end
end

//
genvar i;
// vc_credit_to_return: flag bit per vc to indicate if a vc credit should be returned
generate for (i = 0; i < 13; i=i+1) begin : vc_cred_ret
	assign vc_credit_to_return[i] = |vc_credit[i][8:3];
end
endgenerate

//////////// VC Credits to return counters

// CD VC Credits
generate for (i = 0; i < 2; i=i+1) begin : CD_VCs
	always@(posedge clk) begin
		if(~rst_n) begin
			vc_credit[i] <= 9'b0;
		end
		else if(link_state[0] | link_state[1]) begin
			vc_credit[i] <= CD_LINK_CREDITS;
		end
		else begin
			vc_credit[i] <= vc_credit[i] - ({9{vc_credit_dec[i]}} & 9'd8) + ({9{rx_vc_fifo_pop[i]}} & CD_CREDIT_INC);
		end
	end
end
endgenerate
generate for (i = 2; i < 6; i=i+1) begin : MD_VCs
	always@(posedge clk) begin
		if(~rst_n) begin
			vc_credit[i] <= 9'b0;
		end
		else if(link_state[0] | link_state[1]) begin
			vc_credit[i] <= MD_LINK_CREDITS;
		end
		else begin
			vc_credit[i] <= vc_credit[i] - ({9{vc_credit_dec[i]}} & 9'd8) + ({9{rx_vc_fifo_pop[i]}} & CD_CREDIT_INC);
		end
	end
end
endgenerate
// CO VC Credits
generate for (i = 6; i < 12; i=i+1) begin : CO_VCs
	always@(posedge clk) begin
		if(~rst_n) begin
			vc_credit[i] <= 9'b0;
		end
		else if(link_state[0] | link_state[1]) begin
			vc_credit[i] <= CO_LINK_CREDITS;
		end
		else begin
			vc_credit[i] <= vc_credit[i] - ({9{vc_credit_dec[i]}} & 9'd8) + ({9{rx_vc_fifo_pop[i]}} & CO_CREDIT_INC);
		end
	end
end
endgenerate
// MOC VC Credit
always@(posedge clk) begin
	if(~rst_n) begin
		vc_credit[12] <= 9'b0;
	end
	else if(link_state[0] | link_state[1]) begin
		vc_credit[12] <= MOC_LINK_CREDITS;
	end
	else begin
		vc_credit[12] <= vc_credit[12] - ({9{vc_credit_dec[12]}} & 9'd8) + ({9{rx_vc_fifo_pop[12]}} & MOC_CREDIT_INC);
	end
end


//////////////////////////////////////////////////////////////////////////
/////////////////////////       Replay Memory        /////////////////////
//////////////////////////////////////////////////////////////////////////
assign replay_mem_we    = link_state_sending[2] && !tx_block_out_t.custom_fields[38] && tx_block_out_ready;
assign replay_mem_din   = tx_block_out;
// replay_mem_waddr: whenever we send non IDLe, non Sync blocks we buffer them in the replay buffer,
// only reset the write address when we in initiation states.
//
always@(posedge clk) begin
	if(~rst_n) begin
		replay_mem_waddr <= 8'b0;
	end
	else begin
		if(replay_mem_we) begin
			replay_mem_waddr <= replay_mem_waddr + 1'b1;
		end
		else if(link_state[0] | link_state[1]) begin
			replay_mem_waddr <= 8'b0;
		end
	end
end

////////////////////////////////

assign last_replay_w    = (next_replay_mem_raddr == tx_seq_minus_1);
assign last_replay_sent = last_replay && tx_block_out_ready;
assign retry_ptr        = replay_mem_raddr;
assign replay_mem_re    = link_state[5] && tx_block_out_ready;
//
always@(posedge clk) begin
	if(~rst_n) begin
		replay_mem_raddr <= 8'b0;
		last_replay      <= 1'b0;
	end
	else begin
		replay_mem_raddr <= next_replay_mem_raddr;
		last_replay      <= last_replay_w;
	end
end

always@(*) begin
	if(replay_mem_re) begin
		next_replay_mem_raddr = replay_mem_raddr + 1'b1;
	end
	else if(link_state[4]) begin
		next_replay_mem_raddr = retry_seq;
	end
	else begin
		next_replay_mem_raddr = replay_mem_raddr;
	end
end


// Replay Buffer: Capacity 256 blocks

mem  #( .DATA_WIDTH( $bits(DataBlock_t) ),
        .ADDR_WIDTH(6))
replay_mem
(
    .clk             (clk),

    // Write Port
    .we              (replay_mem_we),
    .waddr           (replay_mem_waddr),
    .din             (replay_mem_din),

    // Read Port
    .raddr           (next_replay_mem_raddr),
    .dout            (replay_mem_block)
);



endmodule
